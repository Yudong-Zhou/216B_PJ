`timescale 1ns / 1ns
module K3_E216_Delta_Y_update_RTL_TB();
reg  clk, rst; 
wire [287:0] dataOut; 
reg [3455:0] dataIn; 
reg [2:0] configIn; 
reg [35:0] controlIn; 
reg [125:0] gcontrolIn; 
reg [31:0] selectedChannel; 
ArrayTop uut(
.clk(clk),
.rst(rst),
.dataOut(dataOut),
.dataIn(dataIn),
.configIn(configIn),
.controlIn(controlIn),
.gControlIn(gcontrolIn)
);
reg [31:0] node_4 = 32'd3;
reg [31:0] node_6 = 32'd3;
reg [31:0] node_7 = 32'd3;
reg [31:0] node_9 = 32'd3;
reg [31:0] node_10 = 32'd3;
always #1 clk = ~clk;
initial begin
rst = 1'b1;
clk = 1'b1;
dataIn = 0;
gcontrolIn = 0;
configIn = 0;
controlIn = 0;
#20
rst = 1'b0;
// Send in configuration bitstream
configIn =3'b010; 
controlIn =36'b000000000000000010000000000000000000; 
#2
configIn =3'b101; 
controlIn =36'b000000000010000000000000000000000000; 
#2
// This is your output channel 
assign selectedChannel =  dataOut[191:160]; 
// Your input IO Config
//000000000000000000000000000000000000000000000000000000000110000000000000000111000000000000000000000000000000
// Your output IO Config
//000000000000000000
// Put together
// Send in IO Configuration 
gcontrolIn =126'b000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000111000000000000000000000000000000; 
// At latency 0 process input node: 10, 9, . 
// At latency 1 process input node: 7, . 
// At latency 2 process input node: . 
// At latency 3 process input node: 6, . 
// At latency 4 process input node: 4, . 
// 40 cycles of constant data to test functionality 
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_4, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9, node_7,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
// alter data to test input latency 
#40
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,   node_10, node_9,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0, node_6,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
dataIn = {
32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0, node_4,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
dataIn = {32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0,32'd0};

end


endmodule
