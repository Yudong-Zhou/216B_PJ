module CADA_InputBuffer (clk, rst, DataIn, DataOut, Sel);
input clk, rst;
input [323:0] Sel; 
input [3455:0] DataIn; 
output [3455:0] DataOut; 
wire [31:0] lin0_0; 
assign lin0_0 = DataIn[3455:3424]; 
wire [31:0] lin0_1; 
CADA_Reg lR0_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin0_0),
.DataOut_1(lin0_1)
);
wire [31:0] lin0_2; 
CADA_Reg lR0_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin0_1),
.DataOut_1(lin0_2)
);
wire [31:0] lin0_3; 
CADA_Reg lR0_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin0_2),
.DataOut_1(lin0_3)
);
wire [31:0] lin0_4; 
CADA_Reg lR0_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin0_3),
.DataOut_1(lin0_4)
);
wire [31:0] lin0_5; 
CADA_Reg lR0_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin0_4),
.DataOut_1(lin0_5)
);
wire [31:0] lout0; 
wire [2:0] sel0; 
HA_6IM lm0(
.sel(sel0),
.DataOut_1(lout0),
.DataIn_1(lin0_0),
.DataIn_2(lin0_1),
.DataIn_3(lin0_2),
.DataIn_4(lin0_3),
.DataIn_5(lin0_4),
.DataIn_6(lin0_5)
);
assign DataOut[3455:3424] = lout0; 
assign sel0 = Sel[323:321]; 
wire [31:0] lin1_0; 
assign lin1_0 = DataIn[3423:3392]; 
wire [31:0] lin1_1; 
CADA_Reg lR1_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin1_0),
.DataOut_1(lin1_1)
);
wire [31:0] lin1_2; 
CADA_Reg lR1_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin1_1),
.DataOut_1(lin1_2)
);
wire [31:0] lin1_3; 
CADA_Reg lR1_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin1_2),
.DataOut_1(lin1_3)
);
wire [31:0] lin1_4; 
CADA_Reg lR1_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin1_3),
.DataOut_1(lin1_4)
);
wire [31:0] lin1_5; 
CADA_Reg lR1_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin1_4),
.DataOut_1(lin1_5)
);
wire [31:0] lout1; 
wire [2:0] sel1; 
HA_6IM lm1(
.sel(sel1),
.DataOut_1(lout1),
.DataIn_1(lin1_0),
.DataIn_2(lin1_1),
.DataIn_3(lin1_2),
.DataIn_4(lin1_3),
.DataIn_5(lin1_4),
.DataIn_6(lin1_5)
);
assign DataOut[3423:3392] = lout1; 
assign sel1 = Sel[320:318]; 
wire [31:0] lin2_0; 
assign lin2_0 = DataIn[3391:3360]; 
wire [31:0] lin2_1; 
CADA_Reg lR2_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin2_0),
.DataOut_1(lin2_1)
);
wire [31:0] lin2_2; 
CADA_Reg lR2_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin2_1),
.DataOut_1(lin2_2)
);
wire [31:0] lin2_3; 
CADA_Reg lR2_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin2_2),
.DataOut_1(lin2_3)
);
wire [31:0] lin2_4; 
CADA_Reg lR2_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin2_3),
.DataOut_1(lin2_4)
);
wire [31:0] lin2_5; 
CADA_Reg lR2_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin2_4),
.DataOut_1(lin2_5)
);
wire [31:0] lout2; 
wire [2:0] sel2; 
HA_6IM lm2(
.sel(sel2),
.DataOut_1(lout2),
.DataIn_1(lin2_0),
.DataIn_2(lin2_1),
.DataIn_3(lin2_2),
.DataIn_4(lin2_3),
.DataIn_5(lin2_4),
.DataIn_6(lin2_5)
);
assign DataOut[3391:3360] = lout2; 
assign sel2 = Sel[317:315]; 
wire [31:0] lin3_0; 
assign lin3_0 = DataIn[3359:3328]; 
wire [31:0] lin3_1; 
CADA_Reg lR3_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin3_0),
.DataOut_1(lin3_1)
);
wire [31:0] lin3_2; 
CADA_Reg lR3_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin3_1),
.DataOut_1(lin3_2)
);
wire [31:0] lin3_3; 
CADA_Reg lR3_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin3_2),
.DataOut_1(lin3_3)
);
wire [31:0] lin3_4; 
CADA_Reg lR3_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin3_3),
.DataOut_1(lin3_4)
);
wire [31:0] lin3_5; 
CADA_Reg lR3_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin3_4),
.DataOut_1(lin3_5)
);
wire [31:0] lout3; 
wire [2:0] sel3; 
HA_6IM lm3(
.sel(sel3),
.DataOut_1(lout3),
.DataIn_1(lin3_0),
.DataIn_2(lin3_1),
.DataIn_3(lin3_2),
.DataIn_4(lin3_3),
.DataIn_5(lin3_4),
.DataIn_6(lin3_5)
);
assign DataOut[3359:3328] = lout3; 
assign sel3 = Sel[314:312]; 
wire [31:0] lin4_0; 
assign lin4_0 = DataIn[3327:3296]; 
wire [31:0] lin4_1; 
CADA_Reg lR4_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin4_0),
.DataOut_1(lin4_1)
);
wire [31:0] lin4_2; 
CADA_Reg lR4_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin4_1),
.DataOut_1(lin4_2)
);
wire [31:0] lin4_3; 
CADA_Reg lR4_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin4_2),
.DataOut_1(lin4_3)
);
wire [31:0] lin4_4; 
CADA_Reg lR4_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin4_3),
.DataOut_1(lin4_4)
);
wire [31:0] lin4_5; 
CADA_Reg lR4_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin4_4),
.DataOut_1(lin4_5)
);
wire [31:0] lout4; 
wire [2:0] sel4; 
HA_6IM lm4(
.sel(sel4),
.DataOut_1(lout4),
.DataIn_1(lin4_0),
.DataIn_2(lin4_1),
.DataIn_3(lin4_2),
.DataIn_4(lin4_3),
.DataIn_5(lin4_4),
.DataIn_6(lin4_5)
);
assign DataOut[3327:3296] = lout4; 
assign sel4 = Sel[311:309]; 
wire [31:0] lin5_0; 
assign lin5_0 = DataIn[3295:3264]; 
wire [31:0] lin5_1; 
CADA_Reg lR5_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin5_0),
.DataOut_1(lin5_1)
);
wire [31:0] lin5_2; 
CADA_Reg lR5_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin5_1),
.DataOut_1(lin5_2)
);
wire [31:0] lin5_3; 
CADA_Reg lR5_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin5_2),
.DataOut_1(lin5_3)
);
wire [31:0] lin5_4; 
CADA_Reg lR5_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin5_3),
.DataOut_1(lin5_4)
);
wire [31:0] lin5_5; 
CADA_Reg lR5_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin5_4),
.DataOut_1(lin5_5)
);
wire [31:0] lout5; 
wire [2:0] sel5; 
HA_6IM lm5(
.sel(sel5),
.DataOut_1(lout5),
.DataIn_1(lin5_0),
.DataIn_2(lin5_1),
.DataIn_3(lin5_2),
.DataIn_4(lin5_3),
.DataIn_5(lin5_4),
.DataIn_6(lin5_5)
);
assign DataOut[3295:3264] = lout5; 
assign sel5 = Sel[308:306]; 
wire [31:0] lin6_0; 
assign lin6_0 = DataIn[3263:3232]; 
wire [31:0] lin6_1; 
CADA_Reg lR6_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin6_0),
.DataOut_1(lin6_1)
);
wire [31:0] lin6_2; 
CADA_Reg lR6_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin6_1),
.DataOut_1(lin6_2)
);
wire [31:0] lin6_3; 
CADA_Reg lR6_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin6_2),
.DataOut_1(lin6_3)
);
wire [31:0] lin6_4; 
CADA_Reg lR6_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin6_3),
.DataOut_1(lin6_4)
);
wire [31:0] lin6_5; 
CADA_Reg lR6_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin6_4),
.DataOut_1(lin6_5)
);
wire [31:0] lout6; 
wire [2:0] sel6; 
HA_6IM lm6(
.sel(sel6),
.DataOut_1(lout6),
.DataIn_1(lin6_0),
.DataIn_2(lin6_1),
.DataIn_3(lin6_2),
.DataIn_4(lin6_3),
.DataIn_5(lin6_4),
.DataIn_6(lin6_5)
);
assign DataOut[3263:3232] = lout6; 
assign sel6 = Sel[305:303]; 
wire [31:0] lin7_0; 
assign lin7_0 = DataIn[3231:3200]; 
wire [31:0] lin7_1; 
CADA_Reg lR7_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin7_0),
.DataOut_1(lin7_1)
);
wire [31:0] lin7_2; 
CADA_Reg lR7_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin7_1),
.DataOut_1(lin7_2)
);
wire [31:0] lin7_3; 
CADA_Reg lR7_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin7_2),
.DataOut_1(lin7_3)
);
wire [31:0] lin7_4; 
CADA_Reg lR7_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin7_3),
.DataOut_1(lin7_4)
);
wire [31:0] lin7_5; 
CADA_Reg lR7_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin7_4),
.DataOut_1(lin7_5)
);
wire [31:0] lout7; 
wire [2:0] sel7; 
HA_6IM lm7(
.sel(sel7),
.DataOut_1(lout7),
.DataIn_1(lin7_0),
.DataIn_2(lin7_1),
.DataIn_3(lin7_2),
.DataIn_4(lin7_3),
.DataIn_5(lin7_4),
.DataIn_6(lin7_5)
);
assign DataOut[3231:3200] = lout7; 
assign sel7 = Sel[302:300]; 
wire [31:0] lin8_0; 
assign lin8_0 = DataIn[3199:3168]; 
wire [31:0] lin8_1; 
CADA_Reg lR8_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin8_0),
.DataOut_1(lin8_1)
);
wire [31:0] lin8_2; 
CADA_Reg lR8_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin8_1),
.DataOut_1(lin8_2)
);
wire [31:0] lin8_3; 
CADA_Reg lR8_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin8_2),
.DataOut_1(lin8_3)
);
wire [31:0] lin8_4; 
CADA_Reg lR8_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin8_3),
.DataOut_1(lin8_4)
);
wire [31:0] lin8_5; 
CADA_Reg lR8_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin8_4),
.DataOut_1(lin8_5)
);
wire [31:0] lout8; 
wire [2:0] sel8; 
HA_6IM lm8(
.sel(sel8),
.DataOut_1(lout8),
.DataIn_1(lin8_0),
.DataIn_2(lin8_1),
.DataIn_3(lin8_2),
.DataIn_4(lin8_3),
.DataIn_5(lin8_4),
.DataIn_6(lin8_5)
);
assign DataOut[3199:3168] = lout8; 
assign sel8 = Sel[299:297]; 
wire [31:0] lin9_0; 
assign lin9_0 = DataIn[3167:3136]; 
wire [31:0] lin9_1; 
CADA_Reg lR9_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin9_0),
.DataOut_1(lin9_1)
);
wire [31:0] lin9_2; 
CADA_Reg lR9_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin9_1),
.DataOut_1(lin9_2)
);
wire [31:0] lin9_3; 
CADA_Reg lR9_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin9_2),
.DataOut_1(lin9_3)
);
wire [31:0] lin9_4; 
CADA_Reg lR9_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin9_3),
.DataOut_1(lin9_4)
);
wire [31:0] lin9_5; 
CADA_Reg lR9_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin9_4),
.DataOut_1(lin9_5)
);
wire [31:0] lout9; 
wire [2:0] sel9; 
HA_6IM lm9(
.sel(sel9),
.DataOut_1(lout9),
.DataIn_1(lin9_0),
.DataIn_2(lin9_1),
.DataIn_3(lin9_2),
.DataIn_4(lin9_3),
.DataIn_5(lin9_4),
.DataIn_6(lin9_5)
);
assign DataOut[3167:3136] = lout9; 
assign sel9 = Sel[296:294]; 
wire [31:0] lin10_0; 
assign lin10_0 = DataIn[3135:3104]; 
wire [31:0] lin10_1; 
CADA_Reg lR10_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin10_0),
.DataOut_1(lin10_1)
);
wire [31:0] lin10_2; 
CADA_Reg lR10_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin10_1),
.DataOut_1(lin10_2)
);
wire [31:0] lin10_3; 
CADA_Reg lR10_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin10_2),
.DataOut_1(lin10_3)
);
wire [31:0] lin10_4; 
CADA_Reg lR10_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin10_3),
.DataOut_1(lin10_4)
);
wire [31:0] lin10_5; 
CADA_Reg lR10_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin10_4),
.DataOut_1(lin10_5)
);
wire [31:0] lout10; 
wire [2:0] sel10; 
HA_6IM lm10(
.sel(sel10),
.DataOut_1(lout10),
.DataIn_1(lin10_0),
.DataIn_2(lin10_1),
.DataIn_3(lin10_2),
.DataIn_4(lin10_3),
.DataIn_5(lin10_4),
.DataIn_6(lin10_5)
);
assign DataOut[3135:3104] = lout10; 
assign sel10 = Sel[293:291]; 
wire [31:0] lin11_0; 
assign lin11_0 = DataIn[3103:3072]; 
wire [31:0] lin11_1; 
CADA_Reg lR11_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin11_0),
.DataOut_1(lin11_1)
);
wire [31:0] lin11_2; 
CADA_Reg lR11_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin11_1),
.DataOut_1(lin11_2)
);
wire [31:0] lin11_3; 
CADA_Reg lR11_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin11_2),
.DataOut_1(lin11_3)
);
wire [31:0] lin11_4; 
CADA_Reg lR11_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin11_3),
.DataOut_1(lin11_4)
);
wire [31:0] lin11_5; 
CADA_Reg lR11_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin11_4),
.DataOut_1(lin11_5)
);
wire [31:0] lout11; 
wire [2:0] sel11; 
HA_6IM lm11(
.sel(sel11),
.DataOut_1(lout11),
.DataIn_1(lin11_0),
.DataIn_2(lin11_1),
.DataIn_3(lin11_2),
.DataIn_4(lin11_3),
.DataIn_5(lin11_4),
.DataIn_6(lin11_5)
);
assign DataOut[3103:3072] = lout11; 
assign sel11 = Sel[290:288]; 
wire [31:0] lin12_0; 
assign lin12_0 = DataIn[3071:3040]; 
wire [31:0] lin12_1; 
CADA_Reg lR12_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin12_0),
.DataOut_1(lin12_1)
);
wire [31:0] lin12_2; 
CADA_Reg lR12_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin12_1),
.DataOut_1(lin12_2)
);
wire [31:0] lin12_3; 
CADA_Reg lR12_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin12_2),
.DataOut_1(lin12_3)
);
wire [31:0] lin12_4; 
CADA_Reg lR12_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin12_3),
.DataOut_1(lin12_4)
);
wire [31:0] lin12_5; 
CADA_Reg lR12_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin12_4),
.DataOut_1(lin12_5)
);
wire [31:0] lout12; 
wire [2:0] sel12; 
HA_6IM lm12(
.sel(sel12),
.DataOut_1(lout12),
.DataIn_1(lin12_0),
.DataIn_2(lin12_1),
.DataIn_3(lin12_2),
.DataIn_4(lin12_3),
.DataIn_5(lin12_4),
.DataIn_6(lin12_5)
);
assign DataOut[3071:3040] = lout12; 
assign sel12 = Sel[287:285]; 
wire [31:0] lin13_0; 
assign lin13_0 = DataIn[3039:3008]; 
wire [31:0] lin13_1; 
CADA_Reg lR13_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin13_0),
.DataOut_1(lin13_1)
);
wire [31:0] lin13_2; 
CADA_Reg lR13_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin13_1),
.DataOut_1(lin13_2)
);
wire [31:0] lin13_3; 
CADA_Reg lR13_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin13_2),
.DataOut_1(lin13_3)
);
wire [31:0] lin13_4; 
CADA_Reg lR13_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin13_3),
.DataOut_1(lin13_4)
);
wire [31:0] lin13_5; 
CADA_Reg lR13_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin13_4),
.DataOut_1(lin13_5)
);
wire [31:0] lout13; 
wire [2:0] sel13; 
HA_6IM lm13(
.sel(sel13),
.DataOut_1(lout13),
.DataIn_1(lin13_0),
.DataIn_2(lin13_1),
.DataIn_3(lin13_2),
.DataIn_4(lin13_3),
.DataIn_5(lin13_4),
.DataIn_6(lin13_5)
);
assign DataOut[3039:3008] = lout13; 
assign sel13 = Sel[284:282]; 
wire [31:0] lin14_0; 
assign lin14_0 = DataIn[3007:2976]; 
wire [31:0] lin14_1; 
CADA_Reg lR14_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin14_0),
.DataOut_1(lin14_1)
);
wire [31:0] lin14_2; 
CADA_Reg lR14_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin14_1),
.DataOut_1(lin14_2)
);
wire [31:0] lin14_3; 
CADA_Reg lR14_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin14_2),
.DataOut_1(lin14_3)
);
wire [31:0] lin14_4; 
CADA_Reg lR14_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin14_3),
.DataOut_1(lin14_4)
);
wire [31:0] lin14_5; 
CADA_Reg lR14_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin14_4),
.DataOut_1(lin14_5)
);
wire [31:0] lout14; 
wire [2:0] sel14; 
HA_6IM lm14(
.sel(sel14),
.DataOut_1(lout14),
.DataIn_1(lin14_0),
.DataIn_2(lin14_1),
.DataIn_3(lin14_2),
.DataIn_4(lin14_3),
.DataIn_5(lin14_4),
.DataIn_6(lin14_5)
);
assign DataOut[3007:2976] = lout14; 
assign sel14 = Sel[281:279]; 
wire [31:0] lin15_0; 
assign lin15_0 = DataIn[2975:2944]; 
wire [31:0] lin15_1; 
CADA_Reg lR15_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin15_0),
.DataOut_1(lin15_1)
);
wire [31:0] lin15_2; 
CADA_Reg lR15_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin15_1),
.DataOut_1(lin15_2)
);
wire [31:0] lin15_3; 
CADA_Reg lR15_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin15_2),
.DataOut_1(lin15_3)
);
wire [31:0] lin15_4; 
CADA_Reg lR15_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin15_3),
.DataOut_1(lin15_4)
);
wire [31:0] lin15_5; 
CADA_Reg lR15_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin15_4),
.DataOut_1(lin15_5)
);
wire [31:0] lout15; 
wire [2:0] sel15; 
HA_6IM lm15(
.sel(sel15),
.DataOut_1(lout15),
.DataIn_1(lin15_0),
.DataIn_2(lin15_1),
.DataIn_3(lin15_2),
.DataIn_4(lin15_3),
.DataIn_5(lin15_4),
.DataIn_6(lin15_5)
);
assign DataOut[2975:2944] = lout15; 
assign sel15 = Sel[278:276]; 
wire [31:0] lin16_0; 
assign lin16_0 = DataIn[2943:2912]; 
wire [31:0] lin16_1; 
CADA_Reg lR16_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin16_0),
.DataOut_1(lin16_1)
);
wire [31:0] lin16_2; 
CADA_Reg lR16_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin16_1),
.DataOut_1(lin16_2)
);
wire [31:0] lin16_3; 
CADA_Reg lR16_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin16_2),
.DataOut_1(lin16_3)
);
wire [31:0] lin16_4; 
CADA_Reg lR16_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin16_3),
.DataOut_1(lin16_4)
);
wire [31:0] lin16_5; 
CADA_Reg lR16_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin16_4),
.DataOut_1(lin16_5)
);
wire [31:0] lout16; 
wire [2:0] sel16; 
HA_6IM lm16(
.sel(sel16),
.DataOut_1(lout16),
.DataIn_1(lin16_0),
.DataIn_2(lin16_1),
.DataIn_3(lin16_2),
.DataIn_4(lin16_3),
.DataIn_5(lin16_4),
.DataIn_6(lin16_5)
);
assign DataOut[2943:2912] = lout16; 
assign sel16 = Sel[275:273]; 
wire [31:0] lin17_0; 
assign lin17_0 = DataIn[2911:2880]; 
wire [31:0] lin17_1; 
CADA_Reg lR17_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin17_0),
.DataOut_1(lin17_1)
);
wire [31:0] lin17_2; 
CADA_Reg lR17_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin17_1),
.DataOut_1(lin17_2)
);
wire [31:0] lin17_3; 
CADA_Reg lR17_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin17_2),
.DataOut_1(lin17_3)
);
wire [31:0] lin17_4; 
CADA_Reg lR17_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin17_3),
.DataOut_1(lin17_4)
);
wire [31:0] lin17_5; 
CADA_Reg lR17_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin17_4),
.DataOut_1(lin17_5)
);
wire [31:0] lout17; 
wire [2:0] sel17; 
HA_6IM lm17(
.sel(sel17),
.DataOut_1(lout17),
.DataIn_1(lin17_0),
.DataIn_2(lin17_1),
.DataIn_3(lin17_2),
.DataIn_4(lin17_3),
.DataIn_5(lin17_4),
.DataIn_6(lin17_5)
);
assign DataOut[2911:2880] = lout17; 
assign sel17 = Sel[272:270]; 
wire [31:0] lin18_0; 
assign lin18_0 = DataIn[2879:2848]; 
wire [31:0] lin18_1; 
CADA_Reg lR18_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin18_0),
.DataOut_1(lin18_1)
);
wire [31:0] lin18_2; 
CADA_Reg lR18_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin18_1),
.DataOut_1(lin18_2)
);
wire [31:0] lin18_3; 
CADA_Reg lR18_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin18_2),
.DataOut_1(lin18_3)
);
wire [31:0] lin18_4; 
CADA_Reg lR18_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin18_3),
.DataOut_1(lin18_4)
);
wire [31:0] lin18_5; 
CADA_Reg lR18_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin18_4),
.DataOut_1(lin18_5)
);
wire [31:0] lout18; 
wire [2:0] sel18; 
HA_6IM lm18(
.sel(sel18),
.DataOut_1(lout18),
.DataIn_1(lin18_0),
.DataIn_2(lin18_1),
.DataIn_3(lin18_2),
.DataIn_4(lin18_3),
.DataIn_5(lin18_4),
.DataIn_6(lin18_5)
);
assign DataOut[2879:2848] = lout18; 
assign sel18 = Sel[269:267]; 
wire [31:0] lin19_0; 
assign lin19_0 = DataIn[2847:2816]; 
wire [31:0] lin19_1; 
CADA_Reg lR19_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin19_0),
.DataOut_1(lin19_1)
);
wire [31:0] lin19_2; 
CADA_Reg lR19_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin19_1),
.DataOut_1(lin19_2)
);
wire [31:0] lin19_3; 
CADA_Reg lR19_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin19_2),
.DataOut_1(lin19_3)
);
wire [31:0] lin19_4; 
CADA_Reg lR19_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin19_3),
.DataOut_1(lin19_4)
);
wire [31:0] lin19_5; 
CADA_Reg lR19_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin19_4),
.DataOut_1(lin19_5)
);
wire [31:0] lout19; 
wire [2:0] sel19; 
HA_6IM lm19(
.sel(sel19),
.DataOut_1(lout19),
.DataIn_1(lin19_0),
.DataIn_2(lin19_1),
.DataIn_3(lin19_2),
.DataIn_4(lin19_3),
.DataIn_5(lin19_4),
.DataIn_6(lin19_5)
);
assign DataOut[2847:2816] = lout19; 
assign sel19 = Sel[266:264]; 
wire [31:0] lin20_0; 
assign lin20_0 = DataIn[2815:2784]; 
wire [31:0] lin20_1; 
CADA_Reg lR20_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin20_0),
.DataOut_1(lin20_1)
);
wire [31:0] lin20_2; 
CADA_Reg lR20_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin20_1),
.DataOut_1(lin20_2)
);
wire [31:0] lin20_3; 
CADA_Reg lR20_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin20_2),
.DataOut_1(lin20_3)
);
wire [31:0] lin20_4; 
CADA_Reg lR20_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin20_3),
.DataOut_1(lin20_4)
);
wire [31:0] lin20_5; 
CADA_Reg lR20_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin20_4),
.DataOut_1(lin20_5)
);
wire [31:0] lout20; 
wire [2:0] sel20; 
HA_6IM lm20(
.sel(sel20),
.DataOut_1(lout20),
.DataIn_1(lin20_0),
.DataIn_2(lin20_1),
.DataIn_3(lin20_2),
.DataIn_4(lin20_3),
.DataIn_5(lin20_4),
.DataIn_6(lin20_5)
);
assign DataOut[2815:2784] = lout20; 
assign sel20 = Sel[263:261]; 
wire [31:0] lin21_0; 
assign lin21_0 = DataIn[2783:2752]; 
wire [31:0] lin21_1; 
CADA_Reg lR21_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin21_0),
.DataOut_1(lin21_1)
);
wire [31:0] lin21_2; 
CADA_Reg lR21_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin21_1),
.DataOut_1(lin21_2)
);
wire [31:0] lin21_3; 
CADA_Reg lR21_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin21_2),
.DataOut_1(lin21_3)
);
wire [31:0] lin21_4; 
CADA_Reg lR21_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin21_3),
.DataOut_1(lin21_4)
);
wire [31:0] lin21_5; 
CADA_Reg lR21_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin21_4),
.DataOut_1(lin21_5)
);
wire [31:0] lout21; 
wire [2:0] sel21; 
HA_6IM lm21(
.sel(sel21),
.DataOut_1(lout21),
.DataIn_1(lin21_0),
.DataIn_2(lin21_1),
.DataIn_3(lin21_2),
.DataIn_4(lin21_3),
.DataIn_5(lin21_4),
.DataIn_6(lin21_5)
);
assign DataOut[2783:2752] = lout21; 
assign sel21 = Sel[260:258]; 
wire [31:0] lin22_0; 
assign lin22_0 = DataIn[2751:2720]; 
wire [31:0] lin22_1; 
CADA_Reg lR22_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin22_0),
.DataOut_1(lin22_1)
);
wire [31:0] lin22_2; 
CADA_Reg lR22_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin22_1),
.DataOut_1(lin22_2)
);
wire [31:0] lin22_3; 
CADA_Reg lR22_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin22_2),
.DataOut_1(lin22_3)
);
wire [31:0] lin22_4; 
CADA_Reg lR22_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin22_3),
.DataOut_1(lin22_4)
);
wire [31:0] lin22_5; 
CADA_Reg lR22_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin22_4),
.DataOut_1(lin22_5)
);
wire [31:0] lout22; 
wire [2:0] sel22; 
HA_6IM lm22(
.sel(sel22),
.DataOut_1(lout22),
.DataIn_1(lin22_0),
.DataIn_2(lin22_1),
.DataIn_3(lin22_2),
.DataIn_4(lin22_3),
.DataIn_5(lin22_4),
.DataIn_6(lin22_5)
);
assign DataOut[2751:2720] = lout22; 
assign sel22 = Sel[257:255]; 
wire [31:0] lin23_0; 
assign lin23_0 = DataIn[2719:2688]; 
wire [31:0] lin23_1; 
CADA_Reg lR23_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin23_0),
.DataOut_1(lin23_1)
);
wire [31:0] lin23_2; 
CADA_Reg lR23_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin23_1),
.DataOut_1(lin23_2)
);
wire [31:0] lin23_3; 
CADA_Reg lR23_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin23_2),
.DataOut_1(lin23_3)
);
wire [31:0] lin23_4; 
CADA_Reg lR23_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin23_3),
.DataOut_1(lin23_4)
);
wire [31:0] lin23_5; 
CADA_Reg lR23_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin23_4),
.DataOut_1(lin23_5)
);
wire [31:0] lout23; 
wire [2:0] sel23; 
HA_6IM lm23(
.sel(sel23),
.DataOut_1(lout23),
.DataIn_1(lin23_0),
.DataIn_2(lin23_1),
.DataIn_3(lin23_2),
.DataIn_4(lin23_3),
.DataIn_5(lin23_4),
.DataIn_6(lin23_5)
);
assign DataOut[2719:2688] = lout23; 
assign sel23 = Sel[254:252]; 
wire [31:0] lin24_0; 
assign lin24_0 = DataIn[2687:2656]; 
wire [31:0] lin24_1; 
CADA_Reg lR24_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin24_0),
.DataOut_1(lin24_1)
);
wire [31:0] lin24_2; 
CADA_Reg lR24_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin24_1),
.DataOut_1(lin24_2)
);
wire [31:0] lin24_3; 
CADA_Reg lR24_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin24_2),
.DataOut_1(lin24_3)
);
wire [31:0] lin24_4; 
CADA_Reg lR24_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin24_3),
.DataOut_1(lin24_4)
);
wire [31:0] lin24_5; 
CADA_Reg lR24_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin24_4),
.DataOut_1(lin24_5)
);
wire [31:0] lout24; 
wire [2:0] sel24; 
HA_6IM lm24(
.sel(sel24),
.DataOut_1(lout24),
.DataIn_1(lin24_0),
.DataIn_2(lin24_1),
.DataIn_3(lin24_2),
.DataIn_4(lin24_3),
.DataIn_5(lin24_4),
.DataIn_6(lin24_5)
);
assign DataOut[2687:2656] = lout24; 
assign sel24 = Sel[251:249]; 
wire [31:0] lin25_0; 
assign lin25_0 = DataIn[2655:2624]; 
wire [31:0] lin25_1; 
CADA_Reg lR25_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin25_0),
.DataOut_1(lin25_1)
);
wire [31:0] lin25_2; 
CADA_Reg lR25_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin25_1),
.DataOut_1(lin25_2)
);
wire [31:0] lin25_3; 
CADA_Reg lR25_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin25_2),
.DataOut_1(lin25_3)
);
wire [31:0] lin25_4; 
CADA_Reg lR25_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin25_3),
.DataOut_1(lin25_4)
);
wire [31:0] lin25_5; 
CADA_Reg lR25_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin25_4),
.DataOut_1(lin25_5)
);
wire [31:0] lout25; 
wire [2:0] sel25; 
HA_6IM lm25(
.sel(sel25),
.DataOut_1(lout25),
.DataIn_1(lin25_0),
.DataIn_2(lin25_1),
.DataIn_3(lin25_2),
.DataIn_4(lin25_3),
.DataIn_5(lin25_4),
.DataIn_6(lin25_5)
);
assign DataOut[2655:2624] = lout25; 
assign sel25 = Sel[248:246]; 
wire [31:0] lin26_0; 
assign lin26_0 = DataIn[2623:2592]; 
wire [31:0] lin26_1; 
CADA_Reg lR26_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin26_0),
.DataOut_1(lin26_1)
);
wire [31:0] lin26_2; 
CADA_Reg lR26_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin26_1),
.DataOut_1(lin26_2)
);
wire [31:0] lin26_3; 
CADA_Reg lR26_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin26_2),
.DataOut_1(lin26_3)
);
wire [31:0] lin26_4; 
CADA_Reg lR26_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin26_3),
.DataOut_1(lin26_4)
);
wire [31:0] lin26_5; 
CADA_Reg lR26_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin26_4),
.DataOut_1(lin26_5)
);
wire [31:0] lout26; 
wire [2:0] sel26; 
HA_6IM lm26(
.sel(sel26),
.DataOut_1(lout26),
.DataIn_1(lin26_0),
.DataIn_2(lin26_1),
.DataIn_3(lin26_2),
.DataIn_4(lin26_3),
.DataIn_5(lin26_4),
.DataIn_6(lin26_5)
);
assign DataOut[2623:2592] = lout26; 
assign sel26 = Sel[245:243]; 
wire [31:0] lin27_0; 
assign lin27_0 = DataIn[2591:2560]; 
wire [31:0] lin27_1; 
CADA_Reg lR27_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin27_0),
.DataOut_1(lin27_1)
);
wire [31:0] lin27_2; 
CADA_Reg lR27_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin27_1),
.DataOut_1(lin27_2)
);
wire [31:0] lin27_3; 
CADA_Reg lR27_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin27_2),
.DataOut_1(lin27_3)
);
wire [31:0] lin27_4; 
CADA_Reg lR27_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin27_3),
.DataOut_1(lin27_4)
);
wire [31:0] lin27_5; 
CADA_Reg lR27_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin27_4),
.DataOut_1(lin27_5)
);
wire [31:0] lout27; 
wire [2:0] sel27; 
HA_6IM lm27(
.sel(sel27),
.DataOut_1(lout27),
.DataIn_1(lin27_0),
.DataIn_2(lin27_1),
.DataIn_3(lin27_2),
.DataIn_4(lin27_3),
.DataIn_5(lin27_4),
.DataIn_6(lin27_5)
);
assign DataOut[2591:2560] = lout27; 
assign sel27 = Sel[242:240]; 
wire [31:0] lin28_0; 
assign lin28_0 = DataIn[2559:2528]; 
wire [31:0] lin28_1; 
CADA_Reg lR28_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin28_0),
.DataOut_1(lin28_1)
);
wire [31:0] lin28_2; 
CADA_Reg lR28_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin28_1),
.DataOut_1(lin28_2)
);
wire [31:0] lin28_3; 
CADA_Reg lR28_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin28_2),
.DataOut_1(lin28_3)
);
wire [31:0] lin28_4; 
CADA_Reg lR28_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin28_3),
.DataOut_1(lin28_4)
);
wire [31:0] lin28_5; 
CADA_Reg lR28_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin28_4),
.DataOut_1(lin28_5)
);
wire [31:0] lout28; 
wire [2:0] sel28; 
HA_6IM lm28(
.sel(sel28),
.DataOut_1(lout28),
.DataIn_1(lin28_0),
.DataIn_2(lin28_1),
.DataIn_3(lin28_2),
.DataIn_4(lin28_3),
.DataIn_5(lin28_4),
.DataIn_6(lin28_5)
);
assign DataOut[2559:2528] = lout28; 
assign sel28 = Sel[239:237]; 
wire [31:0] lin29_0; 
assign lin29_0 = DataIn[2527:2496]; 
wire [31:0] lin29_1; 
CADA_Reg lR29_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin29_0),
.DataOut_1(lin29_1)
);
wire [31:0] lin29_2; 
CADA_Reg lR29_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin29_1),
.DataOut_1(lin29_2)
);
wire [31:0] lin29_3; 
CADA_Reg lR29_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin29_2),
.DataOut_1(lin29_3)
);
wire [31:0] lin29_4; 
CADA_Reg lR29_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin29_3),
.DataOut_1(lin29_4)
);
wire [31:0] lin29_5; 
CADA_Reg lR29_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin29_4),
.DataOut_1(lin29_5)
);
wire [31:0] lout29; 
wire [2:0] sel29; 
HA_6IM lm29(
.sel(sel29),
.DataOut_1(lout29),
.DataIn_1(lin29_0),
.DataIn_2(lin29_1),
.DataIn_3(lin29_2),
.DataIn_4(lin29_3),
.DataIn_5(lin29_4),
.DataIn_6(lin29_5)
);
assign DataOut[2527:2496] = lout29; 
assign sel29 = Sel[236:234]; 
wire [31:0] lin30_0; 
assign lin30_0 = DataIn[2495:2464]; 
wire [31:0] lin30_1; 
CADA_Reg lR30_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin30_0),
.DataOut_1(lin30_1)
);
wire [31:0] lin30_2; 
CADA_Reg lR30_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin30_1),
.DataOut_1(lin30_2)
);
wire [31:0] lin30_3; 
CADA_Reg lR30_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin30_2),
.DataOut_1(lin30_3)
);
wire [31:0] lin30_4; 
CADA_Reg lR30_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin30_3),
.DataOut_1(lin30_4)
);
wire [31:0] lin30_5; 
CADA_Reg lR30_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin30_4),
.DataOut_1(lin30_5)
);
wire [31:0] lout30; 
wire [2:0] sel30; 
HA_6IM lm30(
.sel(sel30),
.DataOut_1(lout30),
.DataIn_1(lin30_0),
.DataIn_2(lin30_1),
.DataIn_3(lin30_2),
.DataIn_4(lin30_3),
.DataIn_5(lin30_4),
.DataIn_6(lin30_5)
);
assign DataOut[2495:2464] = lout30; 
assign sel30 = Sel[233:231]; 
wire [31:0] lin31_0; 
assign lin31_0 = DataIn[2463:2432]; 
wire [31:0] lin31_1; 
CADA_Reg lR31_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin31_0),
.DataOut_1(lin31_1)
);
wire [31:0] lin31_2; 
CADA_Reg lR31_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin31_1),
.DataOut_1(lin31_2)
);
wire [31:0] lin31_3; 
CADA_Reg lR31_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin31_2),
.DataOut_1(lin31_3)
);
wire [31:0] lin31_4; 
CADA_Reg lR31_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin31_3),
.DataOut_1(lin31_4)
);
wire [31:0] lin31_5; 
CADA_Reg lR31_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin31_4),
.DataOut_1(lin31_5)
);
wire [31:0] lout31; 
wire [2:0] sel31; 
HA_6IM lm31(
.sel(sel31),
.DataOut_1(lout31),
.DataIn_1(lin31_0),
.DataIn_2(lin31_1),
.DataIn_3(lin31_2),
.DataIn_4(lin31_3),
.DataIn_5(lin31_4),
.DataIn_6(lin31_5)
);
assign DataOut[2463:2432] = lout31; 
assign sel31 = Sel[230:228]; 
wire [31:0] lin32_0; 
assign lin32_0 = DataIn[2431:2400]; 
wire [31:0] lin32_1; 
CADA_Reg lR32_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin32_0),
.DataOut_1(lin32_1)
);
wire [31:0] lin32_2; 
CADA_Reg lR32_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin32_1),
.DataOut_1(lin32_2)
);
wire [31:0] lin32_3; 
CADA_Reg lR32_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin32_2),
.DataOut_1(lin32_3)
);
wire [31:0] lin32_4; 
CADA_Reg lR32_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin32_3),
.DataOut_1(lin32_4)
);
wire [31:0] lin32_5; 
CADA_Reg lR32_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin32_4),
.DataOut_1(lin32_5)
);
wire [31:0] lout32; 
wire [2:0] sel32; 
HA_6IM lm32(
.sel(sel32),
.DataOut_1(lout32),
.DataIn_1(lin32_0),
.DataIn_2(lin32_1),
.DataIn_3(lin32_2),
.DataIn_4(lin32_3),
.DataIn_5(lin32_4),
.DataIn_6(lin32_5)
);
assign DataOut[2431:2400] = lout32; 
assign sel32 = Sel[227:225]; 
wire [31:0] lin33_0; 
assign lin33_0 = DataIn[2399:2368]; 
wire [31:0] lin33_1; 
CADA_Reg lR33_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin33_0),
.DataOut_1(lin33_1)
);
wire [31:0] lin33_2; 
CADA_Reg lR33_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin33_1),
.DataOut_1(lin33_2)
);
wire [31:0] lin33_3; 
CADA_Reg lR33_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin33_2),
.DataOut_1(lin33_3)
);
wire [31:0] lin33_4; 
CADA_Reg lR33_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin33_3),
.DataOut_1(lin33_4)
);
wire [31:0] lin33_5; 
CADA_Reg lR33_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin33_4),
.DataOut_1(lin33_5)
);
wire [31:0] lout33; 
wire [2:0] sel33; 
HA_6IM lm33(
.sel(sel33),
.DataOut_1(lout33),
.DataIn_1(lin33_0),
.DataIn_2(lin33_1),
.DataIn_3(lin33_2),
.DataIn_4(lin33_3),
.DataIn_5(lin33_4),
.DataIn_6(lin33_5)
);
assign DataOut[2399:2368] = lout33; 
assign sel33 = Sel[224:222]; 
wire [31:0] lin34_0; 
assign lin34_0 = DataIn[2367:2336]; 
wire [31:0] lin34_1; 
CADA_Reg lR34_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin34_0),
.DataOut_1(lin34_1)
);
wire [31:0] lin34_2; 
CADA_Reg lR34_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin34_1),
.DataOut_1(lin34_2)
);
wire [31:0] lin34_3; 
CADA_Reg lR34_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin34_2),
.DataOut_1(lin34_3)
);
wire [31:0] lin34_4; 
CADA_Reg lR34_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin34_3),
.DataOut_1(lin34_4)
);
wire [31:0] lin34_5; 
CADA_Reg lR34_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin34_4),
.DataOut_1(lin34_5)
);
wire [31:0] lout34; 
wire [2:0] sel34; 
HA_6IM lm34(
.sel(sel34),
.DataOut_1(lout34),
.DataIn_1(lin34_0),
.DataIn_2(lin34_1),
.DataIn_3(lin34_2),
.DataIn_4(lin34_3),
.DataIn_5(lin34_4),
.DataIn_6(lin34_5)
);
assign DataOut[2367:2336] = lout34; 
assign sel34 = Sel[221:219]; 
wire [31:0] lin35_0; 
assign lin35_0 = DataIn[2335:2304]; 
wire [31:0] lin35_1; 
CADA_Reg lR35_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin35_0),
.DataOut_1(lin35_1)
);
wire [31:0] lin35_2; 
CADA_Reg lR35_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin35_1),
.DataOut_1(lin35_2)
);
wire [31:0] lin35_3; 
CADA_Reg lR35_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin35_2),
.DataOut_1(lin35_3)
);
wire [31:0] lin35_4; 
CADA_Reg lR35_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin35_3),
.DataOut_1(lin35_4)
);
wire [31:0] lin35_5; 
CADA_Reg lR35_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin35_4),
.DataOut_1(lin35_5)
);
wire [31:0] lout35; 
wire [2:0] sel35; 
HA_6IM lm35(
.sel(sel35),
.DataOut_1(lout35),
.DataIn_1(lin35_0),
.DataIn_2(lin35_1),
.DataIn_3(lin35_2),
.DataIn_4(lin35_3),
.DataIn_5(lin35_4),
.DataIn_6(lin35_5)
);
assign DataOut[2335:2304] = lout35; 
assign sel35 = Sel[218:216]; 
wire [31:0] lin36_0; 
assign lin36_0 = DataIn[2303:2272]; 
wire [31:0] lin36_1; 
CADA_Reg lR36_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin36_0),
.DataOut_1(lin36_1)
);
wire [31:0] lin36_2; 
CADA_Reg lR36_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin36_1),
.DataOut_1(lin36_2)
);
wire [31:0] lin36_3; 
CADA_Reg lR36_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin36_2),
.DataOut_1(lin36_3)
);
wire [31:0] lin36_4; 
CADA_Reg lR36_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin36_3),
.DataOut_1(lin36_4)
);
wire [31:0] lin36_5; 
CADA_Reg lR36_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin36_4),
.DataOut_1(lin36_5)
);
wire [31:0] lout36; 
wire [2:0] sel36; 
HA_6IM lm36(
.sel(sel36),
.DataOut_1(lout36),
.DataIn_1(lin36_0),
.DataIn_2(lin36_1),
.DataIn_3(lin36_2),
.DataIn_4(lin36_3),
.DataIn_5(lin36_4),
.DataIn_6(lin36_5)
);
assign DataOut[2303:2272] = lout36; 
assign sel36 = Sel[215:213]; 
wire [31:0] lin37_0; 
assign lin37_0 = DataIn[2271:2240]; 
wire [31:0] lin37_1; 
CADA_Reg lR37_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin37_0),
.DataOut_1(lin37_1)
);
wire [31:0] lin37_2; 
CADA_Reg lR37_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin37_1),
.DataOut_1(lin37_2)
);
wire [31:0] lin37_3; 
CADA_Reg lR37_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin37_2),
.DataOut_1(lin37_3)
);
wire [31:0] lin37_4; 
CADA_Reg lR37_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin37_3),
.DataOut_1(lin37_4)
);
wire [31:0] lin37_5; 
CADA_Reg lR37_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin37_4),
.DataOut_1(lin37_5)
);
wire [31:0] lout37; 
wire [2:0] sel37; 
HA_6IM lm37(
.sel(sel37),
.DataOut_1(lout37),
.DataIn_1(lin37_0),
.DataIn_2(lin37_1),
.DataIn_3(lin37_2),
.DataIn_4(lin37_3),
.DataIn_5(lin37_4),
.DataIn_6(lin37_5)
);
assign DataOut[2271:2240] = lout37; 
assign sel37 = Sel[212:210]; 
wire [31:0] lin38_0; 
assign lin38_0 = DataIn[2239:2208]; 
wire [31:0] lin38_1; 
CADA_Reg lR38_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin38_0),
.DataOut_1(lin38_1)
);
wire [31:0] lin38_2; 
CADA_Reg lR38_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin38_1),
.DataOut_1(lin38_2)
);
wire [31:0] lin38_3; 
CADA_Reg lR38_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin38_2),
.DataOut_1(lin38_3)
);
wire [31:0] lin38_4; 
CADA_Reg lR38_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin38_3),
.DataOut_1(lin38_4)
);
wire [31:0] lin38_5; 
CADA_Reg lR38_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin38_4),
.DataOut_1(lin38_5)
);
wire [31:0] lout38; 
wire [2:0] sel38; 
HA_6IM lm38(
.sel(sel38),
.DataOut_1(lout38),
.DataIn_1(lin38_0),
.DataIn_2(lin38_1),
.DataIn_3(lin38_2),
.DataIn_4(lin38_3),
.DataIn_5(lin38_4),
.DataIn_6(lin38_5)
);
assign DataOut[2239:2208] = lout38; 
assign sel38 = Sel[209:207]; 
wire [31:0] lin39_0; 
assign lin39_0 = DataIn[2207:2176]; 
wire [31:0] lin39_1; 
CADA_Reg lR39_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin39_0),
.DataOut_1(lin39_1)
);
wire [31:0] lin39_2; 
CADA_Reg lR39_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin39_1),
.DataOut_1(lin39_2)
);
wire [31:0] lin39_3; 
CADA_Reg lR39_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin39_2),
.DataOut_1(lin39_3)
);
wire [31:0] lin39_4; 
CADA_Reg lR39_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin39_3),
.DataOut_1(lin39_4)
);
wire [31:0] lin39_5; 
CADA_Reg lR39_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin39_4),
.DataOut_1(lin39_5)
);
wire [31:0] lout39; 
wire [2:0] sel39; 
HA_6IM lm39(
.sel(sel39),
.DataOut_1(lout39),
.DataIn_1(lin39_0),
.DataIn_2(lin39_1),
.DataIn_3(lin39_2),
.DataIn_4(lin39_3),
.DataIn_5(lin39_4),
.DataIn_6(lin39_5)
);
assign DataOut[2207:2176] = lout39; 
assign sel39 = Sel[206:204]; 
wire [31:0] lin40_0; 
assign lin40_0 = DataIn[2175:2144]; 
wire [31:0] lin40_1; 
CADA_Reg lR40_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin40_0),
.DataOut_1(lin40_1)
);
wire [31:0] lin40_2; 
CADA_Reg lR40_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin40_1),
.DataOut_1(lin40_2)
);
wire [31:0] lin40_3; 
CADA_Reg lR40_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin40_2),
.DataOut_1(lin40_3)
);
wire [31:0] lin40_4; 
CADA_Reg lR40_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin40_3),
.DataOut_1(lin40_4)
);
wire [31:0] lin40_5; 
CADA_Reg lR40_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin40_4),
.DataOut_1(lin40_5)
);
wire [31:0] lout40; 
wire [2:0] sel40; 
HA_6IM lm40(
.sel(sel40),
.DataOut_1(lout40),
.DataIn_1(lin40_0),
.DataIn_2(lin40_1),
.DataIn_3(lin40_2),
.DataIn_4(lin40_3),
.DataIn_5(lin40_4),
.DataIn_6(lin40_5)
);
assign DataOut[2175:2144] = lout40; 
assign sel40 = Sel[203:201]; 
wire [31:0] lin41_0; 
assign lin41_0 = DataIn[2143:2112]; 
wire [31:0] lin41_1; 
CADA_Reg lR41_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin41_0),
.DataOut_1(lin41_1)
);
wire [31:0] lin41_2; 
CADA_Reg lR41_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin41_1),
.DataOut_1(lin41_2)
);
wire [31:0] lin41_3; 
CADA_Reg lR41_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin41_2),
.DataOut_1(lin41_3)
);
wire [31:0] lin41_4; 
CADA_Reg lR41_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin41_3),
.DataOut_1(lin41_4)
);
wire [31:0] lin41_5; 
CADA_Reg lR41_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin41_4),
.DataOut_1(lin41_5)
);
wire [31:0] lout41; 
wire [2:0] sel41; 
HA_6IM lm41(
.sel(sel41),
.DataOut_1(lout41),
.DataIn_1(lin41_0),
.DataIn_2(lin41_1),
.DataIn_3(lin41_2),
.DataIn_4(lin41_3),
.DataIn_5(lin41_4),
.DataIn_6(lin41_5)
);
assign DataOut[2143:2112] = lout41; 
assign sel41 = Sel[200:198]; 
wire [31:0] lin42_0; 
assign lin42_0 = DataIn[2111:2080]; 
wire [31:0] lin42_1; 
CADA_Reg lR42_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin42_0),
.DataOut_1(lin42_1)
);
wire [31:0] lin42_2; 
CADA_Reg lR42_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin42_1),
.DataOut_1(lin42_2)
);
wire [31:0] lin42_3; 
CADA_Reg lR42_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin42_2),
.DataOut_1(lin42_3)
);
wire [31:0] lin42_4; 
CADA_Reg lR42_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin42_3),
.DataOut_1(lin42_4)
);
wire [31:0] lin42_5; 
CADA_Reg lR42_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin42_4),
.DataOut_1(lin42_5)
);
wire [31:0] lout42; 
wire [2:0] sel42; 
HA_6IM lm42(
.sel(sel42),
.DataOut_1(lout42),
.DataIn_1(lin42_0),
.DataIn_2(lin42_1),
.DataIn_3(lin42_2),
.DataIn_4(lin42_3),
.DataIn_5(lin42_4),
.DataIn_6(lin42_5)
);
assign DataOut[2111:2080] = lout42; 
assign sel42 = Sel[197:195]; 
wire [31:0] lin43_0; 
assign lin43_0 = DataIn[2079:2048]; 
wire [31:0] lin43_1; 
CADA_Reg lR43_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin43_0),
.DataOut_1(lin43_1)
);
wire [31:0] lin43_2; 
CADA_Reg lR43_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin43_1),
.DataOut_1(lin43_2)
);
wire [31:0] lin43_3; 
CADA_Reg lR43_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin43_2),
.DataOut_1(lin43_3)
);
wire [31:0] lin43_4; 
CADA_Reg lR43_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin43_3),
.DataOut_1(lin43_4)
);
wire [31:0] lin43_5; 
CADA_Reg lR43_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin43_4),
.DataOut_1(lin43_5)
);
wire [31:0] lout43; 
wire [2:0] sel43; 
HA_6IM lm43(
.sel(sel43),
.DataOut_1(lout43),
.DataIn_1(lin43_0),
.DataIn_2(lin43_1),
.DataIn_3(lin43_2),
.DataIn_4(lin43_3),
.DataIn_5(lin43_4),
.DataIn_6(lin43_5)
);
assign DataOut[2079:2048] = lout43; 
assign sel43 = Sel[194:192]; 
wire [31:0] lin44_0; 
assign lin44_0 = DataIn[2047:2016]; 
wire [31:0] lin44_1; 
CADA_Reg lR44_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin44_0),
.DataOut_1(lin44_1)
);
wire [31:0] lin44_2; 
CADA_Reg lR44_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin44_1),
.DataOut_1(lin44_2)
);
wire [31:0] lin44_3; 
CADA_Reg lR44_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin44_2),
.DataOut_1(lin44_3)
);
wire [31:0] lin44_4; 
CADA_Reg lR44_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin44_3),
.DataOut_1(lin44_4)
);
wire [31:0] lin44_5; 
CADA_Reg lR44_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin44_4),
.DataOut_1(lin44_5)
);
wire [31:0] lout44; 
wire [2:0] sel44; 
HA_6IM lm44(
.sel(sel44),
.DataOut_1(lout44),
.DataIn_1(lin44_0),
.DataIn_2(lin44_1),
.DataIn_3(lin44_2),
.DataIn_4(lin44_3),
.DataIn_5(lin44_4),
.DataIn_6(lin44_5)
);
assign DataOut[2047:2016] = lout44; 
assign sel44 = Sel[191:189]; 
wire [31:0] lin45_0; 
assign lin45_0 = DataIn[2015:1984]; 
wire [31:0] lin45_1; 
CADA_Reg lR45_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin45_0),
.DataOut_1(lin45_1)
);
wire [31:0] lin45_2; 
CADA_Reg lR45_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin45_1),
.DataOut_1(lin45_2)
);
wire [31:0] lin45_3; 
CADA_Reg lR45_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin45_2),
.DataOut_1(lin45_3)
);
wire [31:0] lin45_4; 
CADA_Reg lR45_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin45_3),
.DataOut_1(lin45_4)
);
wire [31:0] lin45_5; 
CADA_Reg lR45_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin45_4),
.DataOut_1(lin45_5)
);
wire [31:0] lout45; 
wire [2:0] sel45; 
HA_6IM lm45(
.sel(sel45),
.DataOut_1(lout45),
.DataIn_1(lin45_0),
.DataIn_2(lin45_1),
.DataIn_3(lin45_2),
.DataIn_4(lin45_3),
.DataIn_5(lin45_4),
.DataIn_6(lin45_5)
);
assign DataOut[2015:1984] = lout45; 
assign sel45 = Sel[188:186]; 
wire [31:0] lin46_0; 
assign lin46_0 = DataIn[1983:1952]; 
wire [31:0] lin46_1; 
CADA_Reg lR46_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin46_0),
.DataOut_1(lin46_1)
);
wire [31:0] lin46_2; 
CADA_Reg lR46_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin46_1),
.DataOut_1(lin46_2)
);
wire [31:0] lin46_3; 
CADA_Reg lR46_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin46_2),
.DataOut_1(lin46_3)
);
wire [31:0] lin46_4; 
CADA_Reg lR46_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin46_3),
.DataOut_1(lin46_4)
);
wire [31:0] lin46_5; 
CADA_Reg lR46_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin46_4),
.DataOut_1(lin46_5)
);
wire [31:0] lout46; 
wire [2:0] sel46; 
HA_6IM lm46(
.sel(sel46),
.DataOut_1(lout46),
.DataIn_1(lin46_0),
.DataIn_2(lin46_1),
.DataIn_3(lin46_2),
.DataIn_4(lin46_3),
.DataIn_5(lin46_4),
.DataIn_6(lin46_5)
);
assign DataOut[1983:1952] = lout46; 
assign sel46 = Sel[185:183]; 
wire [31:0] lin47_0; 
assign lin47_0 = DataIn[1951:1920]; 
wire [31:0] lin47_1; 
CADA_Reg lR47_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin47_0),
.DataOut_1(lin47_1)
);
wire [31:0] lin47_2; 
CADA_Reg lR47_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin47_1),
.DataOut_1(lin47_2)
);
wire [31:0] lin47_3; 
CADA_Reg lR47_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin47_2),
.DataOut_1(lin47_3)
);
wire [31:0] lin47_4; 
CADA_Reg lR47_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin47_3),
.DataOut_1(lin47_4)
);
wire [31:0] lin47_5; 
CADA_Reg lR47_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin47_4),
.DataOut_1(lin47_5)
);
wire [31:0] lout47; 
wire [2:0] sel47; 
HA_6IM lm47(
.sel(sel47),
.DataOut_1(lout47),
.DataIn_1(lin47_0),
.DataIn_2(lin47_1),
.DataIn_3(lin47_2),
.DataIn_4(lin47_3),
.DataIn_5(lin47_4),
.DataIn_6(lin47_5)
);
assign DataOut[1951:1920] = lout47; 
assign sel47 = Sel[182:180]; 
wire [31:0] lin48_0; 
assign lin48_0 = DataIn[1919:1888]; 
wire [31:0] lin48_1; 
CADA_Reg lR48_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin48_0),
.DataOut_1(lin48_1)
);
wire [31:0] lin48_2; 
CADA_Reg lR48_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin48_1),
.DataOut_1(lin48_2)
);
wire [31:0] lin48_3; 
CADA_Reg lR48_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin48_2),
.DataOut_1(lin48_3)
);
wire [31:0] lin48_4; 
CADA_Reg lR48_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin48_3),
.DataOut_1(lin48_4)
);
wire [31:0] lin48_5; 
CADA_Reg lR48_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin48_4),
.DataOut_1(lin48_5)
);
wire [31:0] lout48; 
wire [2:0] sel48; 
HA_6IM lm48(
.sel(sel48),
.DataOut_1(lout48),
.DataIn_1(lin48_0),
.DataIn_2(lin48_1),
.DataIn_3(lin48_2),
.DataIn_4(lin48_3),
.DataIn_5(lin48_4),
.DataIn_6(lin48_5)
);
assign DataOut[1919:1888] = lout48; 
assign sel48 = Sel[179:177]; 
wire [31:0] lin49_0; 
assign lin49_0 = DataIn[1887:1856]; 
wire [31:0] lin49_1; 
CADA_Reg lR49_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin49_0),
.DataOut_1(lin49_1)
);
wire [31:0] lin49_2; 
CADA_Reg lR49_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin49_1),
.DataOut_1(lin49_2)
);
wire [31:0] lin49_3; 
CADA_Reg lR49_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin49_2),
.DataOut_1(lin49_3)
);
wire [31:0] lin49_4; 
CADA_Reg lR49_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin49_3),
.DataOut_1(lin49_4)
);
wire [31:0] lin49_5; 
CADA_Reg lR49_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin49_4),
.DataOut_1(lin49_5)
);
wire [31:0] lout49; 
wire [2:0] sel49; 
HA_6IM lm49(
.sel(sel49),
.DataOut_1(lout49),
.DataIn_1(lin49_0),
.DataIn_2(lin49_1),
.DataIn_3(lin49_2),
.DataIn_4(lin49_3),
.DataIn_5(lin49_4),
.DataIn_6(lin49_5)
);
assign DataOut[1887:1856] = lout49; 
assign sel49 = Sel[176:174]; 
wire [31:0] lin50_0; 
assign lin50_0 = DataIn[1855:1824]; 
wire [31:0] lin50_1; 
CADA_Reg lR50_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin50_0),
.DataOut_1(lin50_1)
);
wire [31:0] lin50_2; 
CADA_Reg lR50_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin50_1),
.DataOut_1(lin50_2)
);
wire [31:0] lin50_3; 
CADA_Reg lR50_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin50_2),
.DataOut_1(lin50_3)
);
wire [31:0] lin50_4; 
CADA_Reg lR50_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin50_3),
.DataOut_1(lin50_4)
);
wire [31:0] lin50_5; 
CADA_Reg lR50_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin50_4),
.DataOut_1(lin50_5)
);
wire [31:0] lout50; 
wire [2:0] sel50; 
HA_6IM lm50(
.sel(sel50),
.DataOut_1(lout50),
.DataIn_1(lin50_0),
.DataIn_2(lin50_1),
.DataIn_3(lin50_2),
.DataIn_4(lin50_3),
.DataIn_5(lin50_4),
.DataIn_6(lin50_5)
);
assign DataOut[1855:1824] = lout50; 
assign sel50 = Sel[173:171]; 
wire [31:0] lin51_0; 
assign lin51_0 = DataIn[1823:1792]; 
wire [31:0] lin51_1; 
CADA_Reg lR51_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin51_0),
.DataOut_1(lin51_1)
);
wire [31:0] lin51_2; 
CADA_Reg lR51_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin51_1),
.DataOut_1(lin51_2)
);
wire [31:0] lin51_3; 
CADA_Reg lR51_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin51_2),
.DataOut_1(lin51_3)
);
wire [31:0] lin51_4; 
CADA_Reg lR51_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin51_3),
.DataOut_1(lin51_4)
);
wire [31:0] lin51_5; 
CADA_Reg lR51_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin51_4),
.DataOut_1(lin51_5)
);
wire [31:0] lout51; 
wire [2:0] sel51; 
HA_6IM lm51(
.sel(sel51),
.DataOut_1(lout51),
.DataIn_1(lin51_0),
.DataIn_2(lin51_1),
.DataIn_3(lin51_2),
.DataIn_4(lin51_3),
.DataIn_5(lin51_4),
.DataIn_6(lin51_5)
);
assign DataOut[1823:1792] = lout51; 
assign sel51 = Sel[170:168]; 
wire [31:0] lin52_0; 
assign lin52_0 = DataIn[1791:1760]; 
wire [31:0] lin52_1; 
CADA_Reg lR52_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin52_0),
.DataOut_1(lin52_1)
);
wire [31:0] lin52_2; 
CADA_Reg lR52_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin52_1),
.DataOut_1(lin52_2)
);
wire [31:0] lin52_3; 
CADA_Reg lR52_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin52_2),
.DataOut_1(lin52_3)
);
wire [31:0] lin52_4; 
CADA_Reg lR52_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin52_3),
.DataOut_1(lin52_4)
);
wire [31:0] lin52_5; 
CADA_Reg lR52_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin52_4),
.DataOut_1(lin52_5)
);
wire [31:0] lout52; 
wire [2:0] sel52; 
HA_6IM lm52(
.sel(sel52),
.DataOut_1(lout52),
.DataIn_1(lin52_0),
.DataIn_2(lin52_1),
.DataIn_3(lin52_2),
.DataIn_4(lin52_3),
.DataIn_5(lin52_4),
.DataIn_6(lin52_5)
);
assign DataOut[1791:1760] = lout52; 
assign sel52 = Sel[167:165]; 
wire [31:0] lin53_0; 
assign lin53_0 = DataIn[1759:1728]; 
wire [31:0] lin53_1; 
CADA_Reg lR53_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin53_0),
.DataOut_1(lin53_1)
);
wire [31:0] lin53_2; 
CADA_Reg lR53_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin53_1),
.DataOut_1(lin53_2)
);
wire [31:0] lin53_3; 
CADA_Reg lR53_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin53_2),
.DataOut_1(lin53_3)
);
wire [31:0] lin53_4; 
CADA_Reg lR53_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin53_3),
.DataOut_1(lin53_4)
);
wire [31:0] lin53_5; 
CADA_Reg lR53_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin53_4),
.DataOut_1(lin53_5)
);
wire [31:0] lout53; 
wire [2:0] sel53; 
HA_6IM lm53(
.sel(sel53),
.DataOut_1(lout53),
.DataIn_1(lin53_0),
.DataIn_2(lin53_1),
.DataIn_3(lin53_2),
.DataIn_4(lin53_3),
.DataIn_5(lin53_4),
.DataIn_6(lin53_5)
);
assign DataOut[1759:1728] = lout53; 
assign sel53 = Sel[164:162]; 
wire [31:0] lin54_0; 
assign lin54_0 = DataIn[1727:1696]; 
wire [31:0] lin54_1; 
CADA_Reg lR54_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin54_0),
.DataOut_1(lin54_1)
);
wire [31:0] lin54_2; 
CADA_Reg lR54_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin54_1),
.DataOut_1(lin54_2)
);
wire [31:0] lin54_3; 
CADA_Reg lR54_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin54_2),
.DataOut_1(lin54_3)
);
wire [31:0] lin54_4; 
CADA_Reg lR54_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin54_3),
.DataOut_1(lin54_4)
);
wire [31:0] lin54_5; 
CADA_Reg lR54_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin54_4),
.DataOut_1(lin54_5)
);
wire [31:0] lout54; 
wire [2:0] sel54; 
HA_6IM lm54(
.sel(sel54),
.DataOut_1(lout54),
.DataIn_1(lin54_0),
.DataIn_2(lin54_1),
.DataIn_3(lin54_2),
.DataIn_4(lin54_3),
.DataIn_5(lin54_4),
.DataIn_6(lin54_5)
);
assign DataOut[1727:1696] = lout54; 
assign sel54 = Sel[161:159]; 
wire [31:0] lin55_0; 
assign lin55_0 = DataIn[1695:1664]; 
wire [31:0] lin55_1; 
CADA_Reg lR55_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin55_0),
.DataOut_1(lin55_1)
);
wire [31:0] lin55_2; 
CADA_Reg lR55_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin55_1),
.DataOut_1(lin55_2)
);
wire [31:0] lin55_3; 
CADA_Reg lR55_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin55_2),
.DataOut_1(lin55_3)
);
wire [31:0] lin55_4; 
CADA_Reg lR55_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin55_3),
.DataOut_1(lin55_4)
);
wire [31:0] lin55_5; 
CADA_Reg lR55_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin55_4),
.DataOut_1(lin55_5)
);
wire [31:0] lout55; 
wire [2:0] sel55; 
HA_6IM lm55(
.sel(sel55),
.DataOut_1(lout55),
.DataIn_1(lin55_0),
.DataIn_2(lin55_1),
.DataIn_3(lin55_2),
.DataIn_4(lin55_3),
.DataIn_5(lin55_4),
.DataIn_6(lin55_5)
);
assign DataOut[1695:1664] = lout55; 
assign sel55 = Sel[158:156]; 
wire [31:0] lin56_0; 
assign lin56_0 = DataIn[1663:1632]; 
wire [31:0] lin56_1; 
CADA_Reg lR56_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin56_0),
.DataOut_1(lin56_1)
);
wire [31:0] lin56_2; 
CADA_Reg lR56_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin56_1),
.DataOut_1(lin56_2)
);
wire [31:0] lin56_3; 
CADA_Reg lR56_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin56_2),
.DataOut_1(lin56_3)
);
wire [31:0] lin56_4; 
CADA_Reg lR56_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin56_3),
.DataOut_1(lin56_4)
);
wire [31:0] lin56_5; 
CADA_Reg lR56_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin56_4),
.DataOut_1(lin56_5)
);
wire [31:0] lout56; 
wire [2:0] sel56; 
HA_6IM lm56(
.sel(sel56),
.DataOut_1(lout56),
.DataIn_1(lin56_0),
.DataIn_2(lin56_1),
.DataIn_3(lin56_2),
.DataIn_4(lin56_3),
.DataIn_5(lin56_4),
.DataIn_6(lin56_5)
);
assign DataOut[1663:1632] = lout56; 
assign sel56 = Sel[155:153]; 
wire [31:0] lin57_0; 
assign lin57_0 = DataIn[1631:1600]; 
wire [31:0] lin57_1; 
CADA_Reg lR57_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin57_0),
.DataOut_1(lin57_1)
);
wire [31:0] lin57_2; 
CADA_Reg lR57_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin57_1),
.DataOut_1(lin57_2)
);
wire [31:0] lin57_3; 
CADA_Reg lR57_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin57_2),
.DataOut_1(lin57_3)
);
wire [31:0] lin57_4; 
CADA_Reg lR57_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin57_3),
.DataOut_1(lin57_4)
);
wire [31:0] lin57_5; 
CADA_Reg lR57_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin57_4),
.DataOut_1(lin57_5)
);
wire [31:0] lout57; 
wire [2:0] sel57; 
HA_6IM lm57(
.sel(sel57),
.DataOut_1(lout57),
.DataIn_1(lin57_0),
.DataIn_2(lin57_1),
.DataIn_3(lin57_2),
.DataIn_4(lin57_3),
.DataIn_5(lin57_4),
.DataIn_6(lin57_5)
);
assign DataOut[1631:1600] = lout57; 
assign sel57 = Sel[152:150]; 
wire [31:0] lin58_0; 
assign lin58_0 = DataIn[1599:1568]; 
wire [31:0] lin58_1; 
CADA_Reg lR58_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin58_0),
.DataOut_1(lin58_1)
);
wire [31:0] lin58_2; 
CADA_Reg lR58_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin58_1),
.DataOut_1(lin58_2)
);
wire [31:0] lin58_3; 
CADA_Reg lR58_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin58_2),
.DataOut_1(lin58_3)
);
wire [31:0] lin58_4; 
CADA_Reg lR58_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin58_3),
.DataOut_1(lin58_4)
);
wire [31:0] lin58_5; 
CADA_Reg lR58_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin58_4),
.DataOut_1(lin58_5)
);
wire [31:0] lout58; 
wire [2:0] sel58; 
HA_6IM lm58(
.sel(sel58),
.DataOut_1(lout58),
.DataIn_1(lin58_0),
.DataIn_2(lin58_1),
.DataIn_3(lin58_2),
.DataIn_4(lin58_3),
.DataIn_5(lin58_4),
.DataIn_6(lin58_5)
);
assign DataOut[1599:1568] = lout58; 
assign sel58 = Sel[149:147]; 
wire [31:0] lin59_0; 
assign lin59_0 = DataIn[1567:1536]; 
wire [31:0] lin59_1; 
CADA_Reg lR59_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin59_0),
.DataOut_1(lin59_1)
);
wire [31:0] lin59_2; 
CADA_Reg lR59_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin59_1),
.DataOut_1(lin59_2)
);
wire [31:0] lin59_3; 
CADA_Reg lR59_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin59_2),
.DataOut_1(lin59_3)
);
wire [31:0] lin59_4; 
CADA_Reg lR59_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin59_3),
.DataOut_1(lin59_4)
);
wire [31:0] lin59_5; 
CADA_Reg lR59_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin59_4),
.DataOut_1(lin59_5)
);
wire [31:0] lout59; 
wire [2:0] sel59; 
HA_6IM lm59(
.sel(sel59),
.DataOut_1(lout59),
.DataIn_1(lin59_0),
.DataIn_2(lin59_1),
.DataIn_3(lin59_2),
.DataIn_4(lin59_3),
.DataIn_5(lin59_4),
.DataIn_6(lin59_5)
);
assign DataOut[1567:1536] = lout59; 
assign sel59 = Sel[146:144]; 
wire [31:0] lin60_0; 
assign lin60_0 = DataIn[1535:1504]; 
wire [31:0] lin60_1; 
CADA_Reg lR60_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin60_0),
.DataOut_1(lin60_1)
);
wire [31:0] lin60_2; 
CADA_Reg lR60_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin60_1),
.DataOut_1(lin60_2)
);
wire [31:0] lin60_3; 
CADA_Reg lR60_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin60_2),
.DataOut_1(lin60_3)
);
wire [31:0] lin60_4; 
CADA_Reg lR60_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin60_3),
.DataOut_1(lin60_4)
);
wire [31:0] lin60_5; 
CADA_Reg lR60_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin60_4),
.DataOut_1(lin60_5)
);
wire [31:0] lout60; 
wire [2:0] sel60; 
HA_6IM lm60(
.sel(sel60),
.DataOut_1(lout60),
.DataIn_1(lin60_0),
.DataIn_2(lin60_1),
.DataIn_3(lin60_2),
.DataIn_4(lin60_3),
.DataIn_5(lin60_4),
.DataIn_6(lin60_5)
);
assign DataOut[1535:1504] = lout60; 
assign sel60 = Sel[143:141]; 
wire [31:0] lin61_0; 
assign lin61_0 = DataIn[1503:1472]; 
wire [31:0] lin61_1; 
CADA_Reg lR61_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin61_0),
.DataOut_1(lin61_1)
);
wire [31:0] lin61_2; 
CADA_Reg lR61_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin61_1),
.DataOut_1(lin61_2)
);
wire [31:0] lin61_3; 
CADA_Reg lR61_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin61_2),
.DataOut_1(lin61_3)
);
wire [31:0] lin61_4; 
CADA_Reg lR61_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin61_3),
.DataOut_1(lin61_4)
);
wire [31:0] lin61_5; 
CADA_Reg lR61_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin61_4),
.DataOut_1(lin61_5)
);
wire [31:0] lout61; 
wire [2:0] sel61; 
HA_6IM lm61(
.sel(sel61),
.DataOut_1(lout61),
.DataIn_1(lin61_0),
.DataIn_2(lin61_1),
.DataIn_3(lin61_2),
.DataIn_4(lin61_3),
.DataIn_5(lin61_4),
.DataIn_6(lin61_5)
);
assign DataOut[1503:1472] = lout61; 
assign sel61 = Sel[140:138]; 
wire [31:0] lin62_0; 
assign lin62_0 = DataIn[1471:1440]; 
wire [31:0] lin62_1; 
CADA_Reg lR62_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin62_0),
.DataOut_1(lin62_1)
);
wire [31:0] lin62_2; 
CADA_Reg lR62_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin62_1),
.DataOut_1(lin62_2)
);
wire [31:0] lin62_3; 
CADA_Reg lR62_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin62_2),
.DataOut_1(lin62_3)
);
wire [31:0] lin62_4; 
CADA_Reg lR62_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin62_3),
.DataOut_1(lin62_4)
);
wire [31:0] lin62_5; 
CADA_Reg lR62_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin62_4),
.DataOut_1(lin62_5)
);
wire [31:0] lout62; 
wire [2:0] sel62; 
HA_6IM lm62(
.sel(sel62),
.DataOut_1(lout62),
.DataIn_1(lin62_0),
.DataIn_2(lin62_1),
.DataIn_3(lin62_2),
.DataIn_4(lin62_3),
.DataIn_5(lin62_4),
.DataIn_6(lin62_5)
);
assign DataOut[1471:1440] = lout62; 
assign sel62 = Sel[137:135]; 
wire [31:0] lin63_0; 
assign lin63_0 = DataIn[1439:1408]; 
wire [31:0] lin63_1; 
CADA_Reg lR63_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin63_0),
.DataOut_1(lin63_1)
);
wire [31:0] lin63_2; 
CADA_Reg lR63_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin63_1),
.DataOut_1(lin63_2)
);
wire [31:0] lin63_3; 
CADA_Reg lR63_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin63_2),
.DataOut_1(lin63_3)
);
wire [31:0] lin63_4; 
CADA_Reg lR63_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin63_3),
.DataOut_1(lin63_4)
);
wire [31:0] lin63_5; 
CADA_Reg lR63_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin63_4),
.DataOut_1(lin63_5)
);
wire [31:0] lout63; 
wire [2:0] sel63; 
HA_6IM lm63(
.sel(sel63),
.DataOut_1(lout63),
.DataIn_1(lin63_0),
.DataIn_2(lin63_1),
.DataIn_3(lin63_2),
.DataIn_4(lin63_3),
.DataIn_5(lin63_4),
.DataIn_6(lin63_5)
);
assign DataOut[1439:1408] = lout63; 
assign sel63 = Sel[134:132]; 
wire [31:0] lin64_0; 
assign lin64_0 = DataIn[1407:1376]; 
wire [31:0] lin64_1; 
CADA_Reg lR64_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin64_0),
.DataOut_1(lin64_1)
);
wire [31:0] lin64_2; 
CADA_Reg lR64_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin64_1),
.DataOut_1(lin64_2)
);
wire [31:0] lin64_3; 
CADA_Reg lR64_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin64_2),
.DataOut_1(lin64_3)
);
wire [31:0] lin64_4; 
CADA_Reg lR64_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin64_3),
.DataOut_1(lin64_4)
);
wire [31:0] lin64_5; 
CADA_Reg lR64_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin64_4),
.DataOut_1(lin64_5)
);
wire [31:0] lout64; 
wire [2:0] sel64; 
HA_6IM lm64(
.sel(sel64),
.DataOut_1(lout64),
.DataIn_1(lin64_0),
.DataIn_2(lin64_1),
.DataIn_3(lin64_2),
.DataIn_4(lin64_3),
.DataIn_5(lin64_4),
.DataIn_6(lin64_5)
);
assign DataOut[1407:1376] = lout64; 
assign sel64 = Sel[131:129]; 
wire [31:0] lin65_0; 
assign lin65_0 = DataIn[1375:1344]; 
wire [31:0] lin65_1; 
CADA_Reg lR65_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin65_0),
.DataOut_1(lin65_1)
);
wire [31:0] lin65_2; 
CADA_Reg lR65_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin65_1),
.DataOut_1(lin65_2)
);
wire [31:0] lin65_3; 
CADA_Reg lR65_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin65_2),
.DataOut_1(lin65_3)
);
wire [31:0] lin65_4; 
CADA_Reg lR65_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin65_3),
.DataOut_1(lin65_4)
);
wire [31:0] lin65_5; 
CADA_Reg lR65_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin65_4),
.DataOut_1(lin65_5)
);
wire [31:0] lout65; 
wire [2:0] sel65; 
HA_6IM lm65(
.sel(sel65),
.DataOut_1(lout65),
.DataIn_1(lin65_0),
.DataIn_2(lin65_1),
.DataIn_3(lin65_2),
.DataIn_4(lin65_3),
.DataIn_5(lin65_4),
.DataIn_6(lin65_5)
);
assign DataOut[1375:1344] = lout65; 
assign sel65 = Sel[128:126]; 
wire [31:0] lin66_0; 
assign lin66_0 = DataIn[1343:1312]; 
wire [31:0] lin66_1; 
CADA_Reg lR66_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin66_0),
.DataOut_1(lin66_1)
);
wire [31:0] lin66_2; 
CADA_Reg lR66_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin66_1),
.DataOut_1(lin66_2)
);
wire [31:0] lin66_3; 
CADA_Reg lR66_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin66_2),
.DataOut_1(lin66_3)
);
wire [31:0] lin66_4; 
CADA_Reg lR66_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin66_3),
.DataOut_1(lin66_4)
);
wire [31:0] lin66_5; 
CADA_Reg lR66_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin66_4),
.DataOut_1(lin66_5)
);
wire [31:0] lout66; 
wire [2:0] sel66; 
HA_6IM lm66(
.sel(sel66),
.DataOut_1(lout66),
.DataIn_1(lin66_0),
.DataIn_2(lin66_1),
.DataIn_3(lin66_2),
.DataIn_4(lin66_3),
.DataIn_5(lin66_4),
.DataIn_6(lin66_5)
);
assign DataOut[1343:1312] = lout66; 
assign sel66 = Sel[125:123]; 
wire [31:0] lin67_0; 
assign lin67_0 = DataIn[1311:1280]; 
wire [31:0] lin67_1; 
CADA_Reg lR67_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin67_0),
.DataOut_1(lin67_1)
);
wire [31:0] lin67_2; 
CADA_Reg lR67_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin67_1),
.DataOut_1(lin67_2)
);
wire [31:0] lin67_3; 
CADA_Reg lR67_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin67_2),
.DataOut_1(lin67_3)
);
wire [31:0] lin67_4; 
CADA_Reg lR67_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin67_3),
.DataOut_1(lin67_4)
);
wire [31:0] lin67_5; 
CADA_Reg lR67_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin67_4),
.DataOut_1(lin67_5)
);
wire [31:0] lout67; 
wire [2:0] sel67; 
HA_6IM lm67(
.sel(sel67),
.DataOut_1(lout67),
.DataIn_1(lin67_0),
.DataIn_2(lin67_1),
.DataIn_3(lin67_2),
.DataIn_4(lin67_3),
.DataIn_5(lin67_4),
.DataIn_6(lin67_5)
);
assign DataOut[1311:1280] = lout67; 
assign sel67 = Sel[122:120]; 
wire [31:0] lin68_0; 
assign lin68_0 = DataIn[1279:1248]; 
wire [31:0] lin68_1; 
CADA_Reg lR68_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin68_0),
.DataOut_1(lin68_1)
);
wire [31:0] lin68_2; 
CADA_Reg lR68_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin68_1),
.DataOut_1(lin68_2)
);
wire [31:0] lin68_3; 
CADA_Reg lR68_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin68_2),
.DataOut_1(lin68_3)
);
wire [31:0] lin68_4; 
CADA_Reg lR68_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin68_3),
.DataOut_1(lin68_4)
);
wire [31:0] lin68_5; 
CADA_Reg lR68_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin68_4),
.DataOut_1(lin68_5)
);
wire [31:0] lout68; 
wire [2:0] sel68; 
HA_6IM lm68(
.sel(sel68),
.DataOut_1(lout68),
.DataIn_1(lin68_0),
.DataIn_2(lin68_1),
.DataIn_3(lin68_2),
.DataIn_4(lin68_3),
.DataIn_5(lin68_4),
.DataIn_6(lin68_5)
);
assign DataOut[1279:1248] = lout68; 
assign sel68 = Sel[119:117]; 
wire [31:0] lin69_0; 
assign lin69_0 = DataIn[1247:1216]; 
wire [31:0] lin69_1; 
CADA_Reg lR69_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin69_0),
.DataOut_1(lin69_1)
);
wire [31:0] lin69_2; 
CADA_Reg lR69_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin69_1),
.DataOut_1(lin69_2)
);
wire [31:0] lin69_3; 
CADA_Reg lR69_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin69_2),
.DataOut_1(lin69_3)
);
wire [31:0] lin69_4; 
CADA_Reg lR69_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin69_3),
.DataOut_1(lin69_4)
);
wire [31:0] lin69_5; 
CADA_Reg lR69_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin69_4),
.DataOut_1(lin69_5)
);
wire [31:0] lout69; 
wire [2:0] sel69; 
HA_6IM lm69(
.sel(sel69),
.DataOut_1(lout69),
.DataIn_1(lin69_0),
.DataIn_2(lin69_1),
.DataIn_3(lin69_2),
.DataIn_4(lin69_3),
.DataIn_5(lin69_4),
.DataIn_6(lin69_5)
);
assign DataOut[1247:1216] = lout69; 
assign sel69 = Sel[116:114]; 
wire [31:0] lin70_0; 
assign lin70_0 = DataIn[1215:1184]; 
wire [31:0] lin70_1; 
CADA_Reg lR70_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin70_0),
.DataOut_1(lin70_1)
);
wire [31:0] lin70_2; 
CADA_Reg lR70_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin70_1),
.DataOut_1(lin70_2)
);
wire [31:0] lin70_3; 
CADA_Reg lR70_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin70_2),
.DataOut_1(lin70_3)
);
wire [31:0] lin70_4; 
CADA_Reg lR70_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin70_3),
.DataOut_1(lin70_4)
);
wire [31:0] lin70_5; 
CADA_Reg lR70_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin70_4),
.DataOut_1(lin70_5)
);
wire [31:0] lout70; 
wire [2:0] sel70; 
HA_6IM lm70(
.sel(sel70),
.DataOut_1(lout70),
.DataIn_1(lin70_0),
.DataIn_2(lin70_1),
.DataIn_3(lin70_2),
.DataIn_4(lin70_3),
.DataIn_5(lin70_4),
.DataIn_6(lin70_5)
);
assign DataOut[1215:1184] = lout70; 
assign sel70 = Sel[113:111]; 
wire [31:0] lin71_0; 
assign lin71_0 = DataIn[1183:1152]; 
wire [31:0] lin71_1; 
CADA_Reg lR71_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin71_0),
.DataOut_1(lin71_1)
);
wire [31:0] lin71_2; 
CADA_Reg lR71_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin71_1),
.DataOut_1(lin71_2)
);
wire [31:0] lin71_3; 
CADA_Reg lR71_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin71_2),
.DataOut_1(lin71_3)
);
wire [31:0] lin71_4; 
CADA_Reg lR71_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin71_3),
.DataOut_1(lin71_4)
);
wire [31:0] lin71_5; 
CADA_Reg lR71_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin71_4),
.DataOut_1(lin71_5)
);
wire [31:0] lout71; 
wire [2:0] sel71; 
HA_6IM lm71(
.sel(sel71),
.DataOut_1(lout71),
.DataIn_1(lin71_0),
.DataIn_2(lin71_1),
.DataIn_3(lin71_2),
.DataIn_4(lin71_3),
.DataIn_5(lin71_4),
.DataIn_6(lin71_5)
);
assign DataOut[1183:1152] = lout71; 
assign sel71 = Sel[110:108]; 
wire [31:0] lin72_0; 
assign lin72_0 = DataIn[1151:1120]; 
wire [31:0] lin72_1; 
CADA_Reg lR72_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin72_0),
.DataOut_1(lin72_1)
);
wire [31:0] lin72_2; 
CADA_Reg lR72_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin72_1),
.DataOut_1(lin72_2)
);
wire [31:0] lin72_3; 
CADA_Reg lR72_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin72_2),
.DataOut_1(lin72_3)
);
wire [31:0] lin72_4; 
CADA_Reg lR72_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin72_3),
.DataOut_1(lin72_4)
);
wire [31:0] lin72_5; 
CADA_Reg lR72_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin72_4),
.DataOut_1(lin72_5)
);
wire [31:0] lout72; 
wire [2:0] sel72; 
HA_6IM lm72(
.sel(sel72),
.DataOut_1(lout72),
.DataIn_1(lin72_0),
.DataIn_2(lin72_1),
.DataIn_3(lin72_2),
.DataIn_4(lin72_3),
.DataIn_5(lin72_4),
.DataIn_6(lin72_5)
);
assign DataOut[1151:1120] = lout72; 
assign sel72 = Sel[107:105]; 
wire [31:0] lin73_0; 
assign lin73_0 = DataIn[1119:1088]; 
wire [31:0] lin73_1; 
CADA_Reg lR73_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin73_0),
.DataOut_1(lin73_1)
);
wire [31:0] lin73_2; 
CADA_Reg lR73_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin73_1),
.DataOut_1(lin73_2)
);
wire [31:0] lin73_3; 
CADA_Reg lR73_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin73_2),
.DataOut_1(lin73_3)
);
wire [31:0] lin73_4; 
CADA_Reg lR73_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin73_3),
.DataOut_1(lin73_4)
);
wire [31:0] lin73_5; 
CADA_Reg lR73_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin73_4),
.DataOut_1(lin73_5)
);
wire [31:0] lout73; 
wire [2:0] sel73; 
HA_6IM lm73(
.sel(sel73),
.DataOut_1(lout73),
.DataIn_1(lin73_0),
.DataIn_2(lin73_1),
.DataIn_3(lin73_2),
.DataIn_4(lin73_3),
.DataIn_5(lin73_4),
.DataIn_6(lin73_5)
);
assign DataOut[1119:1088] = lout73; 
assign sel73 = Sel[104:102]; 
wire [31:0] lin74_0; 
assign lin74_0 = DataIn[1087:1056]; 
wire [31:0] lin74_1; 
CADA_Reg lR74_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin74_0),
.DataOut_1(lin74_1)
);
wire [31:0] lin74_2; 
CADA_Reg lR74_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin74_1),
.DataOut_1(lin74_2)
);
wire [31:0] lin74_3; 
CADA_Reg lR74_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin74_2),
.DataOut_1(lin74_3)
);
wire [31:0] lin74_4; 
CADA_Reg lR74_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin74_3),
.DataOut_1(lin74_4)
);
wire [31:0] lin74_5; 
CADA_Reg lR74_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin74_4),
.DataOut_1(lin74_5)
);
wire [31:0] lout74; 
wire [2:0] sel74; 
HA_6IM lm74(
.sel(sel74),
.DataOut_1(lout74),
.DataIn_1(lin74_0),
.DataIn_2(lin74_1),
.DataIn_3(lin74_2),
.DataIn_4(lin74_3),
.DataIn_5(lin74_4),
.DataIn_6(lin74_5)
);
assign DataOut[1087:1056] = lout74; 
assign sel74 = Sel[101:99]; 
wire [31:0] lin75_0; 
assign lin75_0 = DataIn[1055:1024]; 
wire [31:0] lin75_1; 
CADA_Reg lR75_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin75_0),
.DataOut_1(lin75_1)
);
wire [31:0] lin75_2; 
CADA_Reg lR75_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin75_1),
.DataOut_1(lin75_2)
);
wire [31:0] lin75_3; 
CADA_Reg lR75_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin75_2),
.DataOut_1(lin75_3)
);
wire [31:0] lin75_4; 
CADA_Reg lR75_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin75_3),
.DataOut_1(lin75_4)
);
wire [31:0] lin75_5; 
CADA_Reg lR75_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin75_4),
.DataOut_1(lin75_5)
);
wire [31:0] lout75; 
wire [2:0] sel75; 
HA_6IM lm75(
.sel(sel75),
.DataOut_1(lout75),
.DataIn_1(lin75_0),
.DataIn_2(lin75_1),
.DataIn_3(lin75_2),
.DataIn_4(lin75_3),
.DataIn_5(lin75_4),
.DataIn_6(lin75_5)
);
assign DataOut[1055:1024] = lout75; 
assign sel75 = Sel[98:96]; 
wire [31:0] lin76_0; 
assign lin76_0 = DataIn[1023:992]; 
wire [31:0] lin76_1; 
CADA_Reg lR76_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin76_0),
.DataOut_1(lin76_1)
);
wire [31:0] lin76_2; 
CADA_Reg lR76_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin76_1),
.DataOut_1(lin76_2)
);
wire [31:0] lin76_3; 
CADA_Reg lR76_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin76_2),
.DataOut_1(lin76_3)
);
wire [31:0] lin76_4; 
CADA_Reg lR76_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin76_3),
.DataOut_1(lin76_4)
);
wire [31:0] lin76_5; 
CADA_Reg lR76_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin76_4),
.DataOut_1(lin76_5)
);
wire [31:0] lout76; 
wire [2:0] sel76; 
HA_6IM lm76(
.sel(sel76),
.DataOut_1(lout76),
.DataIn_1(lin76_0),
.DataIn_2(lin76_1),
.DataIn_3(lin76_2),
.DataIn_4(lin76_3),
.DataIn_5(lin76_4),
.DataIn_6(lin76_5)
);
assign DataOut[1023:992] = lout76; 
assign sel76 = Sel[95:93]; 
wire [31:0] lin77_0; 
assign lin77_0 = DataIn[991:960]; 
wire [31:0] lin77_1; 
CADA_Reg lR77_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin77_0),
.DataOut_1(lin77_1)
);
wire [31:0] lin77_2; 
CADA_Reg lR77_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin77_1),
.DataOut_1(lin77_2)
);
wire [31:0] lin77_3; 
CADA_Reg lR77_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin77_2),
.DataOut_1(lin77_3)
);
wire [31:0] lin77_4; 
CADA_Reg lR77_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin77_3),
.DataOut_1(lin77_4)
);
wire [31:0] lin77_5; 
CADA_Reg lR77_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin77_4),
.DataOut_1(lin77_5)
);
wire [31:0] lout77; 
wire [2:0] sel77; 
HA_6IM lm77(
.sel(sel77),
.DataOut_1(lout77),
.DataIn_1(lin77_0),
.DataIn_2(lin77_1),
.DataIn_3(lin77_2),
.DataIn_4(lin77_3),
.DataIn_5(lin77_4),
.DataIn_6(lin77_5)
);
assign DataOut[991:960] = lout77; 
assign sel77 = Sel[92:90]; 
wire [31:0] lin78_0; 
assign lin78_0 = DataIn[959:928]; 
wire [31:0] lin78_1; 
CADA_Reg lR78_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin78_0),
.DataOut_1(lin78_1)
);
wire [31:0] lin78_2; 
CADA_Reg lR78_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin78_1),
.DataOut_1(lin78_2)
);
wire [31:0] lin78_3; 
CADA_Reg lR78_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin78_2),
.DataOut_1(lin78_3)
);
wire [31:0] lin78_4; 
CADA_Reg lR78_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin78_3),
.DataOut_1(lin78_4)
);
wire [31:0] lin78_5; 
CADA_Reg lR78_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin78_4),
.DataOut_1(lin78_5)
);
wire [31:0] lout78; 
wire [2:0] sel78; 
HA_6IM lm78(
.sel(sel78),
.DataOut_1(lout78),
.DataIn_1(lin78_0),
.DataIn_2(lin78_1),
.DataIn_3(lin78_2),
.DataIn_4(lin78_3),
.DataIn_5(lin78_4),
.DataIn_6(lin78_5)
);
assign DataOut[959:928] = lout78; 
assign sel78 = Sel[89:87]; 
wire [31:0] lin79_0; 
assign lin79_0 = DataIn[927:896]; 
wire [31:0] lin79_1; 
CADA_Reg lR79_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin79_0),
.DataOut_1(lin79_1)
);
wire [31:0] lin79_2; 
CADA_Reg lR79_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin79_1),
.DataOut_1(lin79_2)
);
wire [31:0] lin79_3; 
CADA_Reg lR79_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin79_2),
.DataOut_1(lin79_3)
);
wire [31:0] lin79_4; 
CADA_Reg lR79_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin79_3),
.DataOut_1(lin79_4)
);
wire [31:0] lin79_5; 
CADA_Reg lR79_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin79_4),
.DataOut_1(lin79_5)
);
wire [31:0] lout79; 
wire [2:0] sel79; 
HA_6IM lm79(
.sel(sel79),
.DataOut_1(lout79),
.DataIn_1(lin79_0),
.DataIn_2(lin79_1),
.DataIn_3(lin79_2),
.DataIn_4(lin79_3),
.DataIn_5(lin79_4),
.DataIn_6(lin79_5)
);
assign DataOut[927:896] = lout79; 
assign sel79 = Sel[86:84]; 
wire [31:0] lin80_0; 
assign lin80_0 = DataIn[895:864]; 
wire [31:0] lin80_1; 
CADA_Reg lR80_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin80_0),
.DataOut_1(lin80_1)
);
wire [31:0] lin80_2; 
CADA_Reg lR80_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin80_1),
.DataOut_1(lin80_2)
);
wire [31:0] lin80_3; 
CADA_Reg lR80_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin80_2),
.DataOut_1(lin80_3)
);
wire [31:0] lin80_4; 
CADA_Reg lR80_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin80_3),
.DataOut_1(lin80_4)
);
wire [31:0] lin80_5; 
CADA_Reg lR80_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin80_4),
.DataOut_1(lin80_5)
);
wire [31:0] lout80; 
wire [2:0] sel80; 
HA_6IM lm80(
.sel(sel80),
.DataOut_1(lout80),
.DataIn_1(lin80_0),
.DataIn_2(lin80_1),
.DataIn_3(lin80_2),
.DataIn_4(lin80_3),
.DataIn_5(lin80_4),
.DataIn_6(lin80_5)
);
assign DataOut[895:864] = lout80; 
assign sel80 = Sel[83:81]; 
wire [31:0] lin81_0; 
assign lin81_0 = DataIn[863:832]; 
wire [31:0] lin81_1; 
CADA_Reg lR81_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin81_0),
.DataOut_1(lin81_1)
);
wire [31:0] lin81_2; 
CADA_Reg lR81_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin81_1),
.DataOut_1(lin81_2)
);
wire [31:0] lin81_3; 
CADA_Reg lR81_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin81_2),
.DataOut_1(lin81_3)
);
wire [31:0] lin81_4; 
CADA_Reg lR81_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin81_3),
.DataOut_1(lin81_4)
);
wire [31:0] lin81_5; 
CADA_Reg lR81_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin81_4),
.DataOut_1(lin81_5)
);
wire [31:0] lout81; 
wire [2:0] sel81; 
HA_6IM lm81(
.sel(sel81),
.DataOut_1(lout81),
.DataIn_1(lin81_0),
.DataIn_2(lin81_1),
.DataIn_3(lin81_2),
.DataIn_4(lin81_3),
.DataIn_5(lin81_4),
.DataIn_6(lin81_5)
);
assign DataOut[863:832] = lout81; 
assign sel81 = Sel[80:78]; 
wire [31:0] lin82_0; 
assign lin82_0 = DataIn[831:800]; 
wire [31:0] lin82_1; 
CADA_Reg lR82_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin82_0),
.DataOut_1(lin82_1)
);
wire [31:0] lin82_2; 
CADA_Reg lR82_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin82_1),
.DataOut_1(lin82_2)
);
wire [31:0] lin82_3; 
CADA_Reg lR82_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin82_2),
.DataOut_1(lin82_3)
);
wire [31:0] lin82_4; 
CADA_Reg lR82_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin82_3),
.DataOut_1(lin82_4)
);
wire [31:0] lin82_5; 
CADA_Reg lR82_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin82_4),
.DataOut_1(lin82_5)
);
wire [31:0] lout82; 
wire [2:0] sel82; 
HA_6IM lm82(
.sel(sel82),
.DataOut_1(lout82),
.DataIn_1(lin82_0),
.DataIn_2(lin82_1),
.DataIn_3(lin82_2),
.DataIn_4(lin82_3),
.DataIn_5(lin82_4),
.DataIn_6(lin82_5)
);
assign DataOut[831:800] = lout82; 
assign sel82 = Sel[77:75]; 
wire [31:0] lin83_0; 
assign lin83_0 = DataIn[799:768]; 
wire [31:0] lin83_1; 
CADA_Reg lR83_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin83_0),
.DataOut_1(lin83_1)
);
wire [31:0] lin83_2; 
CADA_Reg lR83_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin83_1),
.DataOut_1(lin83_2)
);
wire [31:0] lin83_3; 
CADA_Reg lR83_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin83_2),
.DataOut_1(lin83_3)
);
wire [31:0] lin83_4; 
CADA_Reg lR83_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin83_3),
.DataOut_1(lin83_4)
);
wire [31:0] lin83_5; 
CADA_Reg lR83_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin83_4),
.DataOut_1(lin83_5)
);
wire [31:0] lout83; 
wire [2:0] sel83; 
HA_6IM lm83(
.sel(sel83),
.DataOut_1(lout83),
.DataIn_1(lin83_0),
.DataIn_2(lin83_1),
.DataIn_3(lin83_2),
.DataIn_4(lin83_3),
.DataIn_5(lin83_4),
.DataIn_6(lin83_5)
);
assign DataOut[799:768] = lout83; 
assign sel83 = Sel[74:72]; 
wire [31:0] lin84_0; 
assign lin84_0 = DataIn[767:736]; 
wire [31:0] lin84_1; 
CADA_Reg lR84_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin84_0),
.DataOut_1(lin84_1)
);
wire [31:0] lin84_2; 
CADA_Reg lR84_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin84_1),
.DataOut_1(lin84_2)
);
wire [31:0] lin84_3; 
CADA_Reg lR84_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin84_2),
.DataOut_1(lin84_3)
);
wire [31:0] lin84_4; 
CADA_Reg lR84_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin84_3),
.DataOut_1(lin84_4)
);
wire [31:0] lin84_5; 
CADA_Reg lR84_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin84_4),
.DataOut_1(lin84_5)
);
wire [31:0] lout84; 
wire [2:0] sel84; 
HA_6IM lm84(
.sel(sel84),
.DataOut_1(lout84),
.DataIn_1(lin84_0),
.DataIn_2(lin84_1),
.DataIn_3(lin84_2),
.DataIn_4(lin84_3),
.DataIn_5(lin84_4),
.DataIn_6(lin84_5)
);
assign DataOut[767:736] = lout84; 
assign sel84 = Sel[71:69]; 
wire [31:0] lin85_0; 
assign lin85_0 = DataIn[735:704]; 
wire [31:0] lin85_1; 
CADA_Reg lR85_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin85_0),
.DataOut_1(lin85_1)
);
wire [31:0] lin85_2; 
CADA_Reg lR85_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin85_1),
.DataOut_1(lin85_2)
);
wire [31:0] lin85_3; 
CADA_Reg lR85_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin85_2),
.DataOut_1(lin85_3)
);
wire [31:0] lin85_4; 
CADA_Reg lR85_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin85_3),
.DataOut_1(lin85_4)
);
wire [31:0] lin85_5; 
CADA_Reg lR85_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin85_4),
.DataOut_1(lin85_5)
);
wire [31:0] lout85; 
wire [2:0] sel85; 
HA_6IM lm85(
.sel(sel85),
.DataOut_1(lout85),
.DataIn_1(lin85_0),
.DataIn_2(lin85_1),
.DataIn_3(lin85_2),
.DataIn_4(lin85_3),
.DataIn_5(lin85_4),
.DataIn_6(lin85_5)
);
assign DataOut[735:704] = lout85; 
assign sel85 = Sel[68:66]; 
wire [31:0] lin86_0; 
assign lin86_0 = DataIn[703:672]; 
wire [31:0] lin86_1; 
CADA_Reg lR86_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin86_0),
.DataOut_1(lin86_1)
);
wire [31:0] lin86_2; 
CADA_Reg lR86_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin86_1),
.DataOut_1(lin86_2)
);
wire [31:0] lin86_3; 
CADA_Reg lR86_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin86_2),
.DataOut_1(lin86_3)
);
wire [31:0] lin86_4; 
CADA_Reg lR86_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin86_3),
.DataOut_1(lin86_4)
);
wire [31:0] lin86_5; 
CADA_Reg lR86_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin86_4),
.DataOut_1(lin86_5)
);
wire [31:0] lout86; 
wire [2:0] sel86; 
HA_6IM lm86(
.sel(sel86),
.DataOut_1(lout86),
.DataIn_1(lin86_0),
.DataIn_2(lin86_1),
.DataIn_3(lin86_2),
.DataIn_4(lin86_3),
.DataIn_5(lin86_4),
.DataIn_6(lin86_5)
);
assign DataOut[703:672] = lout86; 
assign sel86 = Sel[65:63]; 
wire [31:0] lin87_0; 
assign lin87_0 = DataIn[671:640]; 
wire [31:0] lin87_1; 
CADA_Reg lR87_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin87_0),
.DataOut_1(lin87_1)
);
wire [31:0] lin87_2; 
CADA_Reg lR87_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin87_1),
.DataOut_1(lin87_2)
);
wire [31:0] lin87_3; 
CADA_Reg lR87_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin87_2),
.DataOut_1(lin87_3)
);
wire [31:0] lin87_4; 
CADA_Reg lR87_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin87_3),
.DataOut_1(lin87_4)
);
wire [31:0] lin87_5; 
CADA_Reg lR87_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin87_4),
.DataOut_1(lin87_5)
);
wire [31:0] lout87; 
wire [2:0] sel87; 
HA_6IM lm87(
.sel(sel87),
.DataOut_1(lout87),
.DataIn_1(lin87_0),
.DataIn_2(lin87_1),
.DataIn_3(lin87_2),
.DataIn_4(lin87_3),
.DataIn_5(lin87_4),
.DataIn_6(lin87_5)
);
assign DataOut[671:640] = lout87; 
assign sel87 = Sel[62:60]; 
wire [31:0] lin88_0; 
assign lin88_0 = DataIn[639:608]; 
wire [31:0] lin88_1; 
CADA_Reg lR88_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin88_0),
.DataOut_1(lin88_1)
);
wire [31:0] lin88_2; 
CADA_Reg lR88_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin88_1),
.DataOut_1(lin88_2)
);
wire [31:0] lin88_3; 
CADA_Reg lR88_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin88_2),
.DataOut_1(lin88_3)
);
wire [31:0] lin88_4; 
CADA_Reg lR88_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin88_3),
.DataOut_1(lin88_4)
);
wire [31:0] lin88_5; 
CADA_Reg lR88_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin88_4),
.DataOut_1(lin88_5)
);
wire [31:0] lout88; 
wire [2:0] sel88; 
HA_6IM lm88(
.sel(sel88),
.DataOut_1(lout88),
.DataIn_1(lin88_0),
.DataIn_2(lin88_1),
.DataIn_3(lin88_2),
.DataIn_4(lin88_3),
.DataIn_5(lin88_4),
.DataIn_6(lin88_5)
);
assign DataOut[639:608] = lout88; 
assign sel88 = Sel[59:57]; 
wire [31:0] lin89_0; 
assign lin89_0 = DataIn[607:576]; 
wire [31:0] lin89_1; 
CADA_Reg lR89_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin89_0),
.DataOut_1(lin89_1)
);
wire [31:0] lin89_2; 
CADA_Reg lR89_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin89_1),
.DataOut_1(lin89_2)
);
wire [31:0] lin89_3; 
CADA_Reg lR89_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin89_2),
.DataOut_1(lin89_3)
);
wire [31:0] lin89_4; 
CADA_Reg lR89_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin89_3),
.DataOut_1(lin89_4)
);
wire [31:0] lin89_5; 
CADA_Reg lR89_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin89_4),
.DataOut_1(lin89_5)
);
wire [31:0] lout89; 
wire [2:0] sel89; 
HA_6IM lm89(
.sel(sel89),
.DataOut_1(lout89),
.DataIn_1(lin89_0),
.DataIn_2(lin89_1),
.DataIn_3(lin89_2),
.DataIn_4(lin89_3),
.DataIn_5(lin89_4),
.DataIn_6(lin89_5)
);
assign DataOut[607:576] = lout89; 
assign sel89 = Sel[56:54]; 
wire [31:0] lin90_0; 
assign lin90_0 = DataIn[575:544]; 
wire [31:0] lin90_1; 
CADA_Reg lR90_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin90_0),
.DataOut_1(lin90_1)
);
wire [31:0] lin90_2; 
CADA_Reg lR90_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin90_1),
.DataOut_1(lin90_2)
);
wire [31:0] lin90_3; 
CADA_Reg lR90_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin90_2),
.DataOut_1(lin90_3)
);
wire [31:0] lin90_4; 
CADA_Reg lR90_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin90_3),
.DataOut_1(lin90_4)
);
wire [31:0] lin90_5; 
CADA_Reg lR90_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin90_4),
.DataOut_1(lin90_5)
);
wire [31:0] lout90; 
wire [2:0] sel90; 
HA_6IM lm90(
.sel(sel90),
.DataOut_1(lout90),
.DataIn_1(lin90_0),
.DataIn_2(lin90_1),
.DataIn_3(lin90_2),
.DataIn_4(lin90_3),
.DataIn_5(lin90_4),
.DataIn_6(lin90_5)
);
assign DataOut[575:544] = lout90; 
assign sel90 = Sel[53:51]; 
wire [31:0] lin91_0; 
assign lin91_0 = DataIn[543:512]; 
wire [31:0] lin91_1; 
CADA_Reg lR91_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin91_0),
.DataOut_1(lin91_1)
);
wire [31:0] lin91_2; 
CADA_Reg lR91_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin91_1),
.DataOut_1(lin91_2)
);
wire [31:0] lin91_3; 
CADA_Reg lR91_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin91_2),
.DataOut_1(lin91_3)
);
wire [31:0] lin91_4; 
CADA_Reg lR91_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin91_3),
.DataOut_1(lin91_4)
);
wire [31:0] lin91_5; 
CADA_Reg lR91_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin91_4),
.DataOut_1(lin91_5)
);
wire [31:0] lout91; 
wire [2:0] sel91; 
HA_6IM lm91(
.sel(sel91),
.DataOut_1(lout91),
.DataIn_1(lin91_0),
.DataIn_2(lin91_1),
.DataIn_3(lin91_2),
.DataIn_4(lin91_3),
.DataIn_5(lin91_4),
.DataIn_6(lin91_5)
);
assign DataOut[543:512] = lout91; 
assign sel91 = Sel[50:48]; 
wire [31:0] lin92_0; 
assign lin92_0 = DataIn[511:480]; 
wire [31:0] lin92_1; 
CADA_Reg lR92_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin92_0),
.DataOut_1(lin92_1)
);
wire [31:0] lin92_2; 
CADA_Reg lR92_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin92_1),
.DataOut_1(lin92_2)
);
wire [31:0] lin92_3; 
CADA_Reg lR92_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin92_2),
.DataOut_1(lin92_3)
);
wire [31:0] lin92_4; 
CADA_Reg lR92_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin92_3),
.DataOut_1(lin92_4)
);
wire [31:0] lin92_5; 
CADA_Reg lR92_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin92_4),
.DataOut_1(lin92_5)
);
wire [31:0] lout92; 
wire [2:0] sel92; 
HA_6IM lm92(
.sel(sel92),
.DataOut_1(lout92),
.DataIn_1(lin92_0),
.DataIn_2(lin92_1),
.DataIn_3(lin92_2),
.DataIn_4(lin92_3),
.DataIn_5(lin92_4),
.DataIn_6(lin92_5)
);
assign DataOut[511:480] = lout92; 
assign sel92 = Sel[47:45]; 
wire [31:0] lin93_0; 
assign lin93_0 = DataIn[479:448]; 
wire [31:0] lin93_1; 
CADA_Reg lR93_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin93_0),
.DataOut_1(lin93_1)
);
wire [31:0] lin93_2; 
CADA_Reg lR93_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin93_1),
.DataOut_1(lin93_2)
);
wire [31:0] lin93_3; 
CADA_Reg lR93_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin93_2),
.DataOut_1(lin93_3)
);
wire [31:0] lin93_4; 
CADA_Reg lR93_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin93_3),
.DataOut_1(lin93_4)
);
wire [31:0] lin93_5; 
CADA_Reg lR93_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin93_4),
.DataOut_1(lin93_5)
);
wire [31:0] lout93; 
wire [2:0] sel93; 
HA_6IM lm93(
.sel(sel93),
.DataOut_1(lout93),
.DataIn_1(lin93_0),
.DataIn_2(lin93_1),
.DataIn_3(lin93_2),
.DataIn_4(lin93_3),
.DataIn_5(lin93_4),
.DataIn_6(lin93_5)
);
assign DataOut[479:448] = lout93; 
assign sel93 = Sel[44:42]; 
wire [31:0] lin94_0; 
assign lin94_0 = DataIn[447:416]; 
wire [31:0] lin94_1; 
CADA_Reg lR94_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin94_0),
.DataOut_1(lin94_1)
);
wire [31:0] lin94_2; 
CADA_Reg lR94_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin94_1),
.DataOut_1(lin94_2)
);
wire [31:0] lin94_3; 
CADA_Reg lR94_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin94_2),
.DataOut_1(lin94_3)
);
wire [31:0] lin94_4; 
CADA_Reg lR94_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin94_3),
.DataOut_1(lin94_4)
);
wire [31:0] lin94_5; 
CADA_Reg lR94_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin94_4),
.DataOut_1(lin94_5)
);
wire [31:0] lout94; 
wire [2:0] sel94; 
HA_6IM lm94(
.sel(sel94),
.DataOut_1(lout94),
.DataIn_1(lin94_0),
.DataIn_2(lin94_1),
.DataIn_3(lin94_2),
.DataIn_4(lin94_3),
.DataIn_5(lin94_4),
.DataIn_6(lin94_5)
);
assign DataOut[447:416] = lout94; 
assign sel94 = Sel[41:39]; 
wire [31:0] lin95_0; 
assign lin95_0 = DataIn[415:384]; 
wire [31:0] lin95_1; 
CADA_Reg lR95_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin95_0),
.DataOut_1(lin95_1)
);
wire [31:0] lin95_2; 
CADA_Reg lR95_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin95_1),
.DataOut_1(lin95_2)
);
wire [31:0] lin95_3; 
CADA_Reg lR95_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin95_2),
.DataOut_1(lin95_3)
);
wire [31:0] lin95_4; 
CADA_Reg lR95_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin95_3),
.DataOut_1(lin95_4)
);
wire [31:0] lin95_5; 
CADA_Reg lR95_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin95_4),
.DataOut_1(lin95_5)
);
wire [31:0] lout95; 
wire [2:0] sel95; 
HA_6IM lm95(
.sel(sel95),
.DataOut_1(lout95),
.DataIn_1(lin95_0),
.DataIn_2(lin95_1),
.DataIn_3(lin95_2),
.DataIn_4(lin95_3),
.DataIn_5(lin95_4),
.DataIn_6(lin95_5)
);
assign DataOut[415:384] = lout95; 
assign sel95 = Sel[38:36]; 
wire [31:0] lin96_0; 
assign lin96_0 = DataIn[383:352]; 
wire [31:0] lin96_1; 
CADA_Reg lR96_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin96_0),
.DataOut_1(lin96_1)
);
wire [31:0] lin96_2; 
CADA_Reg lR96_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin96_1),
.DataOut_1(lin96_2)
);
wire [31:0] lin96_3; 
CADA_Reg lR96_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin96_2),
.DataOut_1(lin96_3)
);
wire [31:0] lin96_4; 
CADA_Reg lR96_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin96_3),
.DataOut_1(lin96_4)
);
wire [31:0] lin96_5; 
CADA_Reg lR96_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin96_4),
.DataOut_1(lin96_5)
);
wire [31:0] lout96; 
wire [2:0] sel96; 
HA_6IM lm96(
.sel(sel96),
.DataOut_1(lout96),
.DataIn_1(lin96_0),
.DataIn_2(lin96_1),
.DataIn_3(lin96_2),
.DataIn_4(lin96_3),
.DataIn_5(lin96_4),
.DataIn_6(lin96_5)
);
assign DataOut[383:352] = lout96; 
assign sel96 = Sel[35:33]; 
wire [31:0] lin97_0; 
assign lin97_0 = DataIn[351:320]; 
wire [31:0] lin97_1; 
CADA_Reg lR97_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin97_0),
.DataOut_1(lin97_1)
);
wire [31:0] lin97_2; 
CADA_Reg lR97_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin97_1),
.DataOut_1(lin97_2)
);
wire [31:0] lin97_3; 
CADA_Reg lR97_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin97_2),
.DataOut_1(lin97_3)
);
wire [31:0] lin97_4; 
CADA_Reg lR97_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin97_3),
.DataOut_1(lin97_4)
);
wire [31:0] lin97_5; 
CADA_Reg lR97_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin97_4),
.DataOut_1(lin97_5)
);
wire [31:0] lout97; 
wire [2:0] sel97; 
HA_6IM lm97(
.sel(sel97),
.DataOut_1(lout97),
.DataIn_1(lin97_0),
.DataIn_2(lin97_1),
.DataIn_3(lin97_2),
.DataIn_4(lin97_3),
.DataIn_5(lin97_4),
.DataIn_6(lin97_5)
);
assign DataOut[351:320] = lout97; 
assign sel97 = Sel[32:30]; 
wire [31:0] lin98_0; 
assign lin98_0 = DataIn[319:288]; 
wire [31:0] lin98_1; 
CADA_Reg lR98_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin98_0),
.DataOut_1(lin98_1)
);
wire [31:0] lin98_2; 
CADA_Reg lR98_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin98_1),
.DataOut_1(lin98_2)
);
wire [31:0] lin98_3; 
CADA_Reg lR98_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin98_2),
.DataOut_1(lin98_3)
);
wire [31:0] lin98_4; 
CADA_Reg lR98_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin98_3),
.DataOut_1(lin98_4)
);
wire [31:0] lin98_5; 
CADA_Reg lR98_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin98_4),
.DataOut_1(lin98_5)
);
wire [31:0] lout98; 
wire [2:0] sel98; 
HA_6IM lm98(
.sel(sel98),
.DataOut_1(lout98),
.DataIn_1(lin98_0),
.DataIn_2(lin98_1),
.DataIn_3(lin98_2),
.DataIn_4(lin98_3),
.DataIn_5(lin98_4),
.DataIn_6(lin98_5)
);
assign DataOut[319:288] = lout98; 
assign sel98 = Sel[29:27]; 
wire [31:0] lin99_0; 
assign lin99_0 = DataIn[287:256]; 
wire [31:0] lin99_1; 
CADA_Reg lR99_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin99_0),
.DataOut_1(lin99_1)
);
wire [31:0] lin99_2; 
CADA_Reg lR99_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin99_1),
.DataOut_1(lin99_2)
);
wire [31:0] lin99_3; 
CADA_Reg lR99_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin99_2),
.DataOut_1(lin99_3)
);
wire [31:0] lin99_4; 
CADA_Reg lR99_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin99_3),
.DataOut_1(lin99_4)
);
wire [31:0] lin99_5; 
CADA_Reg lR99_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin99_4),
.DataOut_1(lin99_5)
);
wire [31:0] lout99; 
wire [2:0] sel99; 
HA_6IM lm99(
.sel(sel99),
.DataOut_1(lout99),
.DataIn_1(lin99_0),
.DataIn_2(lin99_1),
.DataIn_3(lin99_2),
.DataIn_4(lin99_3),
.DataIn_5(lin99_4),
.DataIn_6(lin99_5)
);
assign DataOut[287:256] = lout99; 
assign sel99 = Sel[26:24]; 
wire [31:0] lin100_0; 
assign lin100_0 = DataIn[255:224]; 
wire [31:0] lin100_1; 
CADA_Reg lR100_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin100_0),
.DataOut_1(lin100_1)
);
wire [31:0] lin100_2; 
CADA_Reg lR100_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin100_1),
.DataOut_1(lin100_2)
);
wire [31:0] lin100_3; 
CADA_Reg lR100_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin100_2),
.DataOut_1(lin100_3)
);
wire [31:0] lin100_4; 
CADA_Reg lR100_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin100_3),
.DataOut_1(lin100_4)
);
wire [31:0] lin100_5; 
CADA_Reg lR100_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin100_4),
.DataOut_1(lin100_5)
);
wire [31:0] lout100; 
wire [2:0] sel100; 
HA_6IM lm100(
.sel(sel100),
.DataOut_1(lout100),
.DataIn_1(lin100_0),
.DataIn_2(lin100_1),
.DataIn_3(lin100_2),
.DataIn_4(lin100_3),
.DataIn_5(lin100_4),
.DataIn_6(lin100_5)
);
assign DataOut[255:224] = lout100; 
assign sel100 = Sel[23:21]; 
wire [31:0] lin101_0; 
assign lin101_0 = DataIn[223:192]; 
wire [31:0] lin101_1; 
CADA_Reg lR101_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin101_0),
.DataOut_1(lin101_1)
);
wire [31:0] lin101_2; 
CADA_Reg lR101_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin101_1),
.DataOut_1(lin101_2)
);
wire [31:0] lin101_3; 
CADA_Reg lR101_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin101_2),
.DataOut_1(lin101_3)
);
wire [31:0] lin101_4; 
CADA_Reg lR101_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin101_3),
.DataOut_1(lin101_4)
);
wire [31:0] lin101_5; 
CADA_Reg lR101_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin101_4),
.DataOut_1(lin101_5)
);
wire [31:0] lout101; 
wire [2:0] sel101; 
HA_6IM lm101(
.sel(sel101),
.DataOut_1(lout101),
.DataIn_1(lin101_0),
.DataIn_2(lin101_1),
.DataIn_3(lin101_2),
.DataIn_4(lin101_3),
.DataIn_5(lin101_4),
.DataIn_6(lin101_5)
);
assign DataOut[223:192] = lout101; 
assign sel101 = Sel[20:18]; 
wire [31:0] lin102_0; 
assign lin102_0 = DataIn[191:160]; 
wire [31:0] lin102_1; 
CADA_Reg lR102_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin102_0),
.DataOut_1(lin102_1)
);
wire [31:0] lin102_2; 
CADA_Reg lR102_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin102_1),
.DataOut_1(lin102_2)
);
wire [31:0] lin102_3; 
CADA_Reg lR102_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin102_2),
.DataOut_1(lin102_3)
);
wire [31:0] lin102_4; 
CADA_Reg lR102_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin102_3),
.DataOut_1(lin102_4)
);
wire [31:0] lin102_5; 
CADA_Reg lR102_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin102_4),
.DataOut_1(lin102_5)
);
wire [31:0] lout102; 
wire [2:0] sel102; 
HA_6IM lm102(
.sel(sel102),
.DataOut_1(lout102),
.DataIn_1(lin102_0),
.DataIn_2(lin102_1),
.DataIn_3(lin102_2),
.DataIn_4(lin102_3),
.DataIn_5(lin102_4),
.DataIn_6(lin102_5)
);
assign DataOut[191:160] = lout102; 
assign sel102 = Sel[17:15]; 
wire [31:0] lin103_0; 
assign lin103_0 = DataIn[159:128]; 
wire [31:0] lin103_1; 
CADA_Reg lR103_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin103_0),
.DataOut_1(lin103_1)
);
wire [31:0] lin103_2; 
CADA_Reg lR103_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin103_1),
.DataOut_1(lin103_2)
);
wire [31:0] lin103_3; 
CADA_Reg lR103_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin103_2),
.DataOut_1(lin103_3)
);
wire [31:0] lin103_4; 
CADA_Reg lR103_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin103_3),
.DataOut_1(lin103_4)
);
wire [31:0] lin103_5; 
CADA_Reg lR103_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin103_4),
.DataOut_1(lin103_5)
);
wire [31:0] lout103; 
wire [2:0] sel103; 
HA_6IM lm103(
.sel(sel103),
.DataOut_1(lout103),
.DataIn_1(lin103_0),
.DataIn_2(lin103_1),
.DataIn_3(lin103_2),
.DataIn_4(lin103_3),
.DataIn_5(lin103_4),
.DataIn_6(lin103_5)
);
assign DataOut[159:128] = lout103; 
assign sel103 = Sel[14:12]; 
wire [31:0] lin104_0; 
assign lin104_0 = DataIn[127:96]; 
wire [31:0] lin104_1; 
CADA_Reg lR104_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin104_0),
.DataOut_1(lin104_1)
);
wire [31:0] lin104_2; 
CADA_Reg lR104_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin104_1),
.DataOut_1(lin104_2)
);
wire [31:0] lin104_3; 
CADA_Reg lR104_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin104_2),
.DataOut_1(lin104_3)
);
wire [31:0] lin104_4; 
CADA_Reg lR104_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin104_3),
.DataOut_1(lin104_4)
);
wire [31:0] lin104_5; 
CADA_Reg lR104_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin104_4),
.DataOut_1(lin104_5)
);
wire [31:0] lout104; 
wire [2:0] sel104; 
HA_6IM lm104(
.sel(sel104),
.DataOut_1(lout104),
.DataIn_1(lin104_0),
.DataIn_2(lin104_1),
.DataIn_3(lin104_2),
.DataIn_4(lin104_3),
.DataIn_5(lin104_4),
.DataIn_6(lin104_5)
);
assign DataOut[127:96] = lout104; 
assign sel104 = Sel[11:9]; 
wire [31:0] lin105_0; 
assign lin105_0 = DataIn[95:64]; 
wire [31:0] lin105_1; 
CADA_Reg lR105_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin105_0),
.DataOut_1(lin105_1)
);
wire [31:0] lin105_2; 
CADA_Reg lR105_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin105_1),
.DataOut_1(lin105_2)
);
wire [31:0] lin105_3; 
CADA_Reg lR105_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin105_2),
.DataOut_1(lin105_3)
);
wire [31:0] lin105_4; 
CADA_Reg lR105_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin105_3),
.DataOut_1(lin105_4)
);
wire [31:0] lin105_5; 
CADA_Reg lR105_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin105_4),
.DataOut_1(lin105_5)
);
wire [31:0] lout105; 
wire [2:0] sel105; 
HA_6IM lm105(
.sel(sel105),
.DataOut_1(lout105),
.DataIn_1(lin105_0),
.DataIn_2(lin105_1),
.DataIn_3(lin105_2),
.DataIn_4(lin105_3),
.DataIn_5(lin105_4),
.DataIn_6(lin105_5)
);
assign DataOut[95:64] = lout105; 
assign sel105 = Sel[8:6]; 
wire [31:0] lin106_0; 
assign lin106_0 = DataIn[63:32]; 
wire [31:0] lin106_1; 
CADA_Reg lR106_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin106_0),
.DataOut_1(lin106_1)
);
wire [31:0] lin106_2; 
CADA_Reg lR106_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin106_1),
.DataOut_1(lin106_2)
);
wire [31:0] lin106_3; 
CADA_Reg lR106_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin106_2),
.DataOut_1(lin106_3)
);
wire [31:0] lin106_4; 
CADA_Reg lR106_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin106_3),
.DataOut_1(lin106_4)
);
wire [31:0] lin106_5; 
CADA_Reg lR106_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin106_4),
.DataOut_1(lin106_5)
);
wire [31:0] lout106; 
wire [2:0] sel106; 
HA_6IM lm106(
.sel(sel106),
.DataOut_1(lout106),
.DataIn_1(lin106_0),
.DataIn_2(lin106_1),
.DataIn_3(lin106_2),
.DataIn_4(lin106_3),
.DataIn_5(lin106_4),
.DataIn_6(lin106_5)
);
assign DataOut[63:32] = lout106; 
assign sel106 = Sel[5:3]; 
wire [31:0] lin107_0; 
assign lin107_0 = DataIn[31:0]; 
wire [31:0] lin107_1; 
CADA_Reg lR107_1(
.clk(clk),
.rst(rst),
.DataIn_1(lin107_0),
.DataOut_1(lin107_1)
);
wire [31:0] lin107_2; 
CADA_Reg lR107_2(
.clk(clk),
.rst(rst),
.DataIn_1(lin107_1),
.DataOut_1(lin107_2)
);
wire [31:0] lin107_3; 
CADA_Reg lR107_3(
.clk(clk),
.rst(rst),
.DataIn_1(lin107_2),
.DataOut_1(lin107_3)
);
wire [31:0] lin107_4; 
CADA_Reg lR107_4(
.clk(clk),
.rst(rst),
.DataIn_1(lin107_3),
.DataOut_1(lin107_4)
);
wire [31:0] lin107_5; 
CADA_Reg lR107_5(
.clk(clk),
.rst(rst),
.DataIn_1(lin107_4),
.DataOut_1(lin107_5)
);
wire [31:0] lout107; 
wire [2:0] sel107; 
HA_6IM lm107(
.sel(sel107),
.DataOut_1(lout107),
.DataIn_1(lin107_0),
.DataIn_2(lin107_1),
.DataIn_3(lin107_2),
.DataIn_4(lin107_3),
.DataIn_5(lin107_4),
.DataIn_6(lin107_5)
);
assign DataOut[31:0] = lout107; 
assign sel107 = Sel[2:0]; 
endmodule