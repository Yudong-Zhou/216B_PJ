`timescale 1ns / 1ns
module CADA_Bd_TB();
reg clk, rst;
reg [755:0] count1, count2;
reg [647:0] addrIn1, addrIn2;
reg [107:0] strideIn1, strideIn2;
reg [107:0] writeEnIn1, writeEnIn2, validIn1, validIn2;
reg [557:0] IOConfig;
reg [3455:0] dataIn;
wire [3455:0] dataOut;
reg [38:0] IdataIn;
wire [38:0] IdataOut;
reg [4:0] IaddrIn1, IaddrIn2;
reg [0:0] IstrideIn1, IstrideIn2;
reg IwriteEnIn1, IvalidIn1, IwriteEnIn2, IvalidIn2;
reg [7:0] Icount1, Icount2;
reg [2:0] configIn; 
reg [35:0] controlIn; 
reg [125:0] gcontrolIn;
reg [431:0] mOutConfig;
reg [31:0] selectedChannel1;
reg [31:0] selectedChannel2;
reg [31:0] selectedChannel3;
CADA_Bd_wrapper uut(
.clk(clk),
.rst(rst),
.IOConfig(IOConfig),
.IaddrIn1(IaddrIn1),
.IaddrIn2(IaddrIn2),
.Icount1(Icount1),
.Icount2(Icount2),
.IdataIn(IdataIn),
.IdataOut(IdataOut),
.IstrideIn1(IstrideIn1),
.IstrideIn2(IstrideIn2),
.IvalidIn1(IvalidIn1),
.IvalidIn2(IvalidIn2),
.IwriteEnIn1(IwriteEnIn1),
.IwriteEnIn2(IwriteEnIn2),
.addrIn1(addrIn1),
.addrIn2(addrIn2),
.count1(count1),
.count2(count2),
.dataIn(dataIn),
.dataOut(dataOut),
.strideIn1(strideIn1),
.strideIn2(strideIn2),
.validIn1(validIn1),
.validIn2(validIn2),
.writeEnIn1(writeEnIn1),
.writeEnIn2(writeEnIn2)
);
reg [31:0] node_4 = 32'd3;
reg [31:0] node_5 = 32'd3;
reg [31:0] node_7 = 32'd3;
reg [31:0] node_8 = 32'd3;
always #1 clk = ~clk;
initial begin
rst = 1'b1;
clk = 1'b1;
dataIn = 0;
addrIn1 = 0;
addrIn2 = 0;
count1 = 0;
count2 = 0;
strideIn1 = 0;
strideIn2 = 0;
writeEnIn1 = 0;
writeEnIn2 = 0;
validIn1 = 0;
validIn2 = 0;
IdataIn = 0;
IaddrIn1 = 0;
IaddrIn2 = 0;
Icount1 = 0;
Icount2 = 0;
IstrideIn1 = 0;
IstrideIn2 = 0;
IwriteEnIn1 = 0;
IwriteEnIn2 = 0;
IvalidIn1 = 0;
IvalidIn2 = 0;
#10
rst = 1'b0;
#10
IaddrIn1 = 0;
Icount1 = 2;
IstrideIn1 = 1;
IwriteEnIn1 = 1;
IvalidIn1 = 1;
// Store configuration bitstream
configIn =3'b000; 
controlIn =36'b000000000000000000001000000000000000; 
IdataIn = {configIn, controlIn}; 
#2
IvalidIn1 = 0;
configIn =3'b101; 
controlIn =36'b000000000000001000000000000000000000; 
IdataIn = {configIn, controlIn}; 
#2
IvalidIn1 = 0;
// Load configuration bitstream and distribute
IaddrIn2 = 0;
Icount2 = 2;
IstrideIn2 = 1;
IwriteEnIn2 = 0;
IvalidIn2 = 1;
#2
IvalidIn2 = 0;
#4
// Your input IO Config
//000000000000000000000000000000000000000000000100000000000000000111000000000000000000000000000000000000000000
// Your output IO Config
//000000001000000000
// Put together
gcontrolIn =126'b000000001000000000000000000000000000000000000000000000000000000100000000000000000111000000000000000000000000000000000000000000; 
// Now let's try to figure out memory network configuration
// When we need to get data from external source (store data into ram), we use this configuration
mOutConfig =432'b100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001; 
// Send in IO Configuration 
IOConfig = {mOutConfig, gcontrolIn}; 
// Let's configure data ram to start reading from external datain port 
addrIn1 = {6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0};
count1 = {7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4};
strideIn1 = {1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1};
writeEnIn1 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
validIn1 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
// At latency 0 process input node: 8, 7, . 
// At latency 1 process input node: 5, . 
// At latency 2 process input node: . 
// At latency 3 process input node: 4, . 
dataIn = {
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,   node_8, node_7,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
validIn1 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
dataIn = {
32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0, node_5,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0};
#2
validIn1 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
dataIn = {
32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0};
#2
validIn1 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
dataIn = {
32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,   node_4,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  
32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0,  32'd0,32'd0,32'd0};
#2
validIn1 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
#2
// Now that data is in ram, let's distribute them to array
// This time, data output is store back to ram, so we need new memory network configuration
// This memory network configuration is choosen because: 
// We are routing output to memory0 which is the input memory for input0 at x=0 , y=0;
// We are routing output to memory1 which is the input memory for input1 at x=0 , y=0;
// We are routing output to memory3 which is the input memory for input0 at x=1 , y=0;
// This is consistent with selectedChannel1,2,3 
mOutConfig =432'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000100; 
IOConfig = {mOutConfig, gcontrolIn}; 
addrIn2 = {6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0};
count2 = {7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4};
strideIn2 = {1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1};
writeEnIn2 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
validIn2 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
// Here we always pull valid to 0 in the next cycle. And we wait for output to reach output memory 
#2
validIn2 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
#16
// Ok, let's store the data at the exact right moment
addrIn1 = {6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0};
count1 = {7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4};
strideIn1 = {1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1};
writeEnIn1 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
validIn1 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
#2
validIn1 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
#20
addrIn2 = {6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0,6'd0};
count2 = {7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4,7'd4};
strideIn2 = {1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1,1'd1};
writeEnIn2 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
validIn2 = {1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1};
#2
validIn2 = {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0};
#6
selectedChannel1 =  dataOut[31:0]; 
selectedChannel2 =  dataOut[63:32]; 
selectedChannel3 =  dataOut[127:96]; 

end


endmodule
