`timescale 1ns / 1ns 
module CGRATop (clk, rst, startAddr1, count1, count2, stride1, WEn1, valid1, startAddr2, stride2, WEn2, valid2, IOConfig, globalDataIn, globalDataOut, IglobalDataIn, IglobalDataOut, IstartAddr1, Istride1, IWEn1, Ivalid1, IstartAddr2, Istride2, IWEn2, Ivalid2,mWEn1, mWEn2, mDataToMem, mDataFromMem, mAddr1, mEn1, mAddr2, mEn2, mIWEn1, mIWEn2, Icount1, Icount2, mIDataFromMem, mIDataToMem, mIAddr1, mIEn1, mIAddr2, mIEn2); 
input clk, rst;
input [755:0] count1, count2;
input [647:0] startAddr1, startAddr2;
input [107:0] stride1, stride2;
input [107:0] WEn1, valid1, WEn2, valid2;
input [557:0] IOConfig;
input [3455:0] globalDataIn;
output [3455:0] globalDataOut;
input [38:0] IglobalDataIn;
output [38:0] IglobalDataOut;
input [4:0] IstartAddr1, IstartAddr2;
input [0:0] Istride1, Istride2;
input IWEn1, Ivalid1, IWEn2, Ivalid2;
input [3455:0] mDataFromMem;
output [3455:0] mDataToMem;
output [107:0] mWEn1, mEn1, mWEn2, mEn2;
output [647:0] mAddr1, mAddr2;
input [38:0] mIDataFromMem;
output [38:0] mIDataToMem;
input [7:0] Icount1, Icount2;
output mIWEn1, mIEn1, mIWEn2, mIEn2;
output [4:0] mIAddr1, mIAddr2;
wire [431:0] mOutConfigW;


//Compute Module Instantiation 
wire [3455:0] dataInW;
wire [287:0] dataOutW;
wire [2:0] configInW;
wire [35:0] controlInW;
wire [125:0] gControlInW;
wire [38:0] totalConfigInW;
assign configInW = totalConfigInW[38:36];
assign controlInW = totalConfigInW[35:0];
ArrayTop computeArray(
.clk(clk),
.rst(rst),
.dataOut(dataOutW),
.dataIn(dataInW),
.configIn(configInW),
.controlIn(controlInW),
.gControlIn(gControlInW));


//Mem Control Instantiation 
wire MEMC0_valid_ctx1;
wire MEMC0_valid_ctx2;
wire [31:0] MEMC0_data_from_Core;
wire [31:0] MEMC0_data_to_Core;
wire [5:0] MEMC0_addr_out_ctx1;
wire MEMC0_write_en_ctx1;
wire MEMC0_write_mem_en_ctx1;
wire MEMC0_mem_en_ctx1;
wire [5:0] MEMC0_start_addr_ctx1;
wire [0:0] MEMC0_stride_ctx1;
wire [5:0] MEMC0_addr_out_ctx2;
wire MEMC0_write_en_ctx2;
wire MEMC0_write_mem_en_ctx2;
wire MEMC0_mem_en_ctx2;
wire [5:0] MEMC0_start_addr_ctx2;
wire [0:0] MEMC0_stride_ctx2;
wire [31:0] MEMC0_data_in_ctx1;
wire [31:0] MEMC0_data_in_ctx2;
wire [31:0] MEMC0_data_out_ctx1;
wire [31:0] MEMC0_data_out_ctx2;
wire [63:0] MEMC0_burst_count_ctx1;
wire [63:0] MEMC0_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC0(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC0_data_from_Core),
.data_to_Core(MEMC0_data_to_Core),
.valid_ctx1(MEMC0_valid_ctx1),
.addr_out_ctx1(MEMC0_addr_out_ctx1),
.write_en_ctx1(MEMC0_write_en_ctx1),
.start_addr_ctx1(MEMC0_start_addr_ctx1),
.stride_ctx1(MEMC0_stride_ctx1),
.burst_count_ctx1(MEMC0_burst_count_ctx1),
.valid_ctx2(MEMC0_valid_ctx2),
.addr_out_ctx2(MEMC0_addr_out_ctx2),
.write_en_ctx2(MEMC0_write_en_ctx2),
.start_addr_ctx2(MEMC0_start_addr_ctx2),
.stride_ctx2(MEMC0_stride_ctx2),
.burst_count_ctx2(MEMC0_burst_count_ctx2),
.data_in_ctx1(MEMC0_data_in_ctx1),
.data_in_ctx2(MEMC0_data_in_ctx2),
.data_out_ctx1(MEMC0_data_out_ctx1),
.data_out_ctx2(MEMC0_data_out_ctx2),
.write_mem_en_ctx1(MEMC0_write_mem_en_ctx1),
.mem_en_ctx1(MEMC0_mem_en_ctx1),.write_mem_en_ctx2(MEMC0_write_mem_en_ctx2),
.mem_en_ctx2(MEMC0_mem_en_ctx2));

defparam MEMC0.DATA_WIDTH = 32;
defparam MEMC0.ADDR_WIDTH = 6;
defparam MEMC0.STRIDE_WIDTH = 1;
wire MEMC1_valid_ctx1;
wire MEMC1_valid_ctx2;
wire [31:0] MEMC1_data_from_Core;
wire [31:0] MEMC1_data_to_Core;
wire [5:0] MEMC1_addr_out_ctx1;
wire MEMC1_write_en_ctx1;
wire MEMC1_write_mem_en_ctx1;
wire MEMC1_mem_en_ctx1;
wire [5:0] MEMC1_start_addr_ctx1;
wire [0:0] MEMC1_stride_ctx1;
wire [5:0] MEMC1_addr_out_ctx2;
wire MEMC1_write_en_ctx2;
wire MEMC1_write_mem_en_ctx2;
wire MEMC1_mem_en_ctx2;
wire [5:0] MEMC1_start_addr_ctx2;
wire [0:0] MEMC1_stride_ctx2;
wire [31:0] MEMC1_data_in_ctx1;
wire [31:0] MEMC1_data_in_ctx2;
wire [31:0] MEMC1_data_out_ctx1;
wire [31:0] MEMC1_data_out_ctx2;
wire [63:0] MEMC1_burst_count_ctx1;
wire [63:0] MEMC1_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC1(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC1_data_from_Core),
.data_to_Core(MEMC1_data_to_Core),
.valid_ctx1(MEMC1_valid_ctx1),
.addr_out_ctx1(MEMC1_addr_out_ctx1),
.write_en_ctx1(MEMC1_write_en_ctx1),
.start_addr_ctx1(MEMC1_start_addr_ctx1),
.stride_ctx1(MEMC1_stride_ctx1),
.burst_count_ctx1(MEMC1_burst_count_ctx1),
.valid_ctx2(MEMC1_valid_ctx2),
.addr_out_ctx2(MEMC1_addr_out_ctx2),
.write_en_ctx2(MEMC1_write_en_ctx2),
.start_addr_ctx2(MEMC1_start_addr_ctx2),
.stride_ctx2(MEMC1_stride_ctx2),
.burst_count_ctx2(MEMC1_burst_count_ctx2),
.data_in_ctx1(MEMC1_data_in_ctx1),
.data_in_ctx2(MEMC1_data_in_ctx2),
.data_out_ctx1(MEMC1_data_out_ctx1),
.data_out_ctx2(MEMC1_data_out_ctx2),
.write_mem_en_ctx1(MEMC1_write_mem_en_ctx1),
.mem_en_ctx1(MEMC1_mem_en_ctx1),.write_mem_en_ctx2(MEMC1_write_mem_en_ctx2),
.mem_en_ctx2(MEMC1_mem_en_ctx2));

defparam MEMC1.DATA_WIDTH = 32;
defparam MEMC1.ADDR_WIDTH = 6;
defparam MEMC1.STRIDE_WIDTH = 1;
wire MEMC2_valid_ctx1;
wire MEMC2_valid_ctx2;
wire [31:0] MEMC2_data_from_Core;
wire [31:0] MEMC2_data_to_Core;
wire [5:0] MEMC2_addr_out_ctx1;
wire MEMC2_write_en_ctx1;
wire MEMC2_write_mem_en_ctx1;
wire MEMC2_mem_en_ctx1;
wire [5:0] MEMC2_start_addr_ctx1;
wire [0:0] MEMC2_stride_ctx1;
wire [5:0] MEMC2_addr_out_ctx2;
wire MEMC2_write_en_ctx2;
wire MEMC2_write_mem_en_ctx2;
wire MEMC2_mem_en_ctx2;
wire [5:0] MEMC2_start_addr_ctx2;
wire [0:0] MEMC2_stride_ctx2;
wire [31:0] MEMC2_data_in_ctx1;
wire [31:0] MEMC2_data_in_ctx2;
wire [31:0] MEMC2_data_out_ctx1;
wire [31:0] MEMC2_data_out_ctx2;
wire [63:0] MEMC2_burst_count_ctx1;
wire [63:0] MEMC2_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC2(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC2_data_from_Core),
.data_to_Core(MEMC2_data_to_Core),
.valid_ctx1(MEMC2_valid_ctx1),
.addr_out_ctx1(MEMC2_addr_out_ctx1),
.write_en_ctx1(MEMC2_write_en_ctx1),
.start_addr_ctx1(MEMC2_start_addr_ctx1),
.stride_ctx1(MEMC2_stride_ctx1),
.burst_count_ctx1(MEMC2_burst_count_ctx1),
.valid_ctx2(MEMC2_valid_ctx2),
.addr_out_ctx2(MEMC2_addr_out_ctx2),
.write_en_ctx2(MEMC2_write_en_ctx2),
.start_addr_ctx2(MEMC2_start_addr_ctx2),
.stride_ctx2(MEMC2_stride_ctx2),
.burst_count_ctx2(MEMC2_burst_count_ctx2),
.data_in_ctx1(MEMC2_data_in_ctx1),
.data_in_ctx2(MEMC2_data_in_ctx2),
.data_out_ctx1(MEMC2_data_out_ctx1),
.data_out_ctx2(MEMC2_data_out_ctx2),
.write_mem_en_ctx1(MEMC2_write_mem_en_ctx1),
.mem_en_ctx1(MEMC2_mem_en_ctx1),.write_mem_en_ctx2(MEMC2_write_mem_en_ctx2),
.mem_en_ctx2(MEMC2_mem_en_ctx2));

defparam MEMC2.DATA_WIDTH = 32;
defparam MEMC2.ADDR_WIDTH = 6;
defparam MEMC2.STRIDE_WIDTH = 1;
wire MEMC3_valid_ctx1;
wire MEMC3_valid_ctx2;
wire [31:0] MEMC3_data_from_Core;
wire [31:0] MEMC3_data_to_Core;
wire [5:0] MEMC3_addr_out_ctx1;
wire MEMC3_write_en_ctx1;
wire MEMC3_write_mem_en_ctx1;
wire MEMC3_mem_en_ctx1;
wire [5:0] MEMC3_start_addr_ctx1;
wire [0:0] MEMC3_stride_ctx1;
wire [5:0] MEMC3_addr_out_ctx2;
wire MEMC3_write_en_ctx2;
wire MEMC3_write_mem_en_ctx2;
wire MEMC3_mem_en_ctx2;
wire [5:0] MEMC3_start_addr_ctx2;
wire [0:0] MEMC3_stride_ctx2;
wire [31:0] MEMC3_data_in_ctx1;
wire [31:0] MEMC3_data_in_ctx2;
wire [31:0] MEMC3_data_out_ctx1;
wire [31:0] MEMC3_data_out_ctx2;
wire [63:0] MEMC3_burst_count_ctx1;
wire [63:0] MEMC3_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC3(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC3_data_from_Core),
.data_to_Core(MEMC3_data_to_Core),
.valid_ctx1(MEMC3_valid_ctx1),
.addr_out_ctx1(MEMC3_addr_out_ctx1),
.write_en_ctx1(MEMC3_write_en_ctx1),
.start_addr_ctx1(MEMC3_start_addr_ctx1),
.stride_ctx1(MEMC3_stride_ctx1),
.burst_count_ctx1(MEMC3_burst_count_ctx1),
.valid_ctx2(MEMC3_valid_ctx2),
.addr_out_ctx2(MEMC3_addr_out_ctx2),
.write_en_ctx2(MEMC3_write_en_ctx2),
.start_addr_ctx2(MEMC3_start_addr_ctx2),
.stride_ctx2(MEMC3_stride_ctx2),
.burst_count_ctx2(MEMC3_burst_count_ctx2),
.data_in_ctx1(MEMC3_data_in_ctx1),
.data_in_ctx2(MEMC3_data_in_ctx2),
.data_out_ctx1(MEMC3_data_out_ctx1),
.data_out_ctx2(MEMC3_data_out_ctx2),
.write_mem_en_ctx1(MEMC3_write_mem_en_ctx1),
.mem_en_ctx1(MEMC3_mem_en_ctx1),.write_mem_en_ctx2(MEMC3_write_mem_en_ctx2),
.mem_en_ctx2(MEMC3_mem_en_ctx2));

defparam MEMC3.DATA_WIDTH = 32;
defparam MEMC3.ADDR_WIDTH = 6;
defparam MEMC3.STRIDE_WIDTH = 1;
wire MEMC4_valid_ctx1;
wire MEMC4_valid_ctx2;
wire [31:0] MEMC4_data_from_Core;
wire [31:0] MEMC4_data_to_Core;
wire [5:0] MEMC4_addr_out_ctx1;
wire MEMC4_write_en_ctx1;
wire MEMC4_write_mem_en_ctx1;
wire MEMC4_mem_en_ctx1;
wire [5:0] MEMC4_start_addr_ctx1;
wire [0:0] MEMC4_stride_ctx1;
wire [5:0] MEMC4_addr_out_ctx2;
wire MEMC4_write_en_ctx2;
wire MEMC4_write_mem_en_ctx2;
wire MEMC4_mem_en_ctx2;
wire [5:0] MEMC4_start_addr_ctx2;
wire [0:0] MEMC4_stride_ctx2;
wire [31:0] MEMC4_data_in_ctx1;
wire [31:0] MEMC4_data_in_ctx2;
wire [31:0] MEMC4_data_out_ctx1;
wire [31:0] MEMC4_data_out_ctx2;
wire [63:0] MEMC4_burst_count_ctx1;
wire [63:0] MEMC4_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC4(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC4_data_from_Core),
.data_to_Core(MEMC4_data_to_Core),
.valid_ctx1(MEMC4_valid_ctx1),
.addr_out_ctx1(MEMC4_addr_out_ctx1),
.write_en_ctx1(MEMC4_write_en_ctx1),
.start_addr_ctx1(MEMC4_start_addr_ctx1),
.stride_ctx1(MEMC4_stride_ctx1),
.burst_count_ctx1(MEMC4_burst_count_ctx1),
.valid_ctx2(MEMC4_valid_ctx2),
.addr_out_ctx2(MEMC4_addr_out_ctx2),
.write_en_ctx2(MEMC4_write_en_ctx2),
.start_addr_ctx2(MEMC4_start_addr_ctx2),
.stride_ctx2(MEMC4_stride_ctx2),
.burst_count_ctx2(MEMC4_burst_count_ctx2),
.data_in_ctx1(MEMC4_data_in_ctx1),
.data_in_ctx2(MEMC4_data_in_ctx2),
.data_out_ctx1(MEMC4_data_out_ctx1),
.data_out_ctx2(MEMC4_data_out_ctx2),
.write_mem_en_ctx1(MEMC4_write_mem_en_ctx1),
.mem_en_ctx1(MEMC4_mem_en_ctx1),.write_mem_en_ctx2(MEMC4_write_mem_en_ctx2),
.mem_en_ctx2(MEMC4_mem_en_ctx2));

defparam MEMC4.DATA_WIDTH = 32;
defparam MEMC4.ADDR_WIDTH = 6;
defparam MEMC4.STRIDE_WIDTH = 1;
wire MEMC5_valid_ctx1;
wire MEMC5_valid_ctx2;
wire [31:0] MEMC5_data_from_Core;
wire [31:0] MEMC5_data_to_Core;
wire [5:0] MEMC5_addr_out_ctx1;
wire MEMC5_write_en_ctx1;
wire MEMC5_write_mem_en_ctx1;
wire MEMC5_mem_en_ctx1;
wire [5:0] MEMC5_start_addr_ctx1;
wire [0:0] MEMC5_stride_ctx1;
wire [5:0] MEMC5_addr_out_ctx2;
wire MEMC5_write_en_ctx2;
wire MEMC5_write_mem_en_ctx2;
wire MEMC5_mem_en_ctx2;
wire [5:0] MEMC5_start_addr_ctx2;
wire [0:0] MEMC5_stride_ctx2;
wire [31:0] MEMC5_data_in_ctx1;
wire [31:0] MEMC5_data_in_ctx2;
wire [31:0] MEMC5_data_out_ctx1;
wire [31:0] MEMC5_data_out_ctx2;
wire [63:0] MEMC5_burst_count_ctx1;
wire [63:0] MEMC5_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC5(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC5_data_from_Core),
.data_to_Core(MEMC5_data_to_Core),
.valid_ctx1(MEMC5_valid_ctx1),
.addr_out_ctx1(MEMC5_addr_out_ctx1),
.write_en_ctx1(MEMC5_write_en_ctx1),
.start_addr_ctx1(MEMC5_start_addr_ctx1),
.stride_ctx1(MEMC5_stride_ctx1),
.burst_count_ctx1(MEMC5_burst_count_ctx1),
.valid_ctx2(MEMC5_valid_ctx2),
.addr_out_ctx2(MEMC5_addr_out_ctx2),
.write_en_ctx2(MEMC5_write_en_ctx2),
.start_addr_ctx2(MEMC5_start_addr_ctx2),
.stride_ctx2(MEMC5_stride_ctx2),
.burst_count_ctx2(MEMC5_burst_count_ctx2),
.data_in_ctx1(MEMC5_data_in_ctx1),
.data_in_ctx2(MEMC5_data_in_ctx2),
.data_out_ctx1(MEMC5_data_out_ctx1),
.data_out_ctx2(MEMC5_data_out_ctx2),
.write_mem_en_ctx1(MEMC5_write_mem_en_ctx1),
.mem_en_ctx1(MEMC5_mem_en_ctx1),.write_mem_en_ctx2(MEMC5_write_mem_en_ctx2),
.mem_en_ctx2(MEMC5_mem_en_ctx2));

defparam MEMC5.DATA_WIDTH = 32;
defparam MEMC5.ADDR_WIDTH = 6;
defparam MEMC5.STRIDE_WIDTH = 1;
wire MEMC6_valid_ctx1;
wire MEMC6_valid_ctx2;
wire [31:0] MEMC6_data_from_Core;
wire [31:0] MEMC6_data_to_Core;
wire [5:0] MEMC6_addr_out_ctx1;
wire MEMC6_write_en_ctx1;
wire MEMC6_write_mem_en_ctx1;
wire MEMC6_mem_en_ctx1;
wire [5:0] MEMC6_start_addr_ctx1;
wire [0:0] MEMC6_stride_ctx1;
wire [5:0] MEMC6_addr_out_ctx2;
wire MEMC6_write_en_ctx2;
wire MEMC6_write_mem_en_ctx2;
wire MEMC6_mem_en_ctx2;
wire [5:0] MEMC6_start_addr_ctx2;
wire [0:0] MEMC6_stride_ctx2;
wire [31:0] MEMC6_data_in_ctx1;
wire [31:0] MEMC6_data_in_ctx2;
wire [31:0] MEMC6_data_out_ctx1;
wire [31:0] MEMC6_data_out_ctx2;
wire [63:0] MEMC6_burst_count_ctx1;
wire [63:0] MEMC6_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC6(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC6_data_from_Core),
.data_to_Core(MEMC6_data_to_Core),
.valid_ctx1(MEMC6_valid_ctx1),
.addr_out_ctx1(MEMC6_addr_out_ctx1),
.write_en_ctx1(MEMC6_write_en_ctx1),
.start_addr_ctx1(MEMC6_start_addr_ctx1),
.stride_ctx1(MEMC6_stride_ctx1),
.burst_count_ctx1(MEMC6_burst_count_ctx1),
.valid_ctx2(MEMC6_valid_ctx2),
.addr_out_ctx2(MEMC6_addr_out_ctx2),
.write_en_ctx2(MEMC6_write_en_ctx2),
.start_addr_ctx2(MEMC6_start_addr_ctx2),
.stride_ctx2(MEMC6_stride_ctx2),
.burst_count_ctx2(MEMC6_burst_count_ctx2),
.data_in_ctx1(MEMC6_data_in_ctx1),
.data_in_ctx2(MEMC6_data_in_ctx2),
.data_out_ctx1(MEMC6_data_out_ctx1),
.data_out_ctx2(MEMC6_data_out_ctx2),
.write_mem_en_ctx1(MEMC6_write_mem_en_ctx1),
.mem_en_ctx1(MEMC6_mem_en_ctx1),.write_mem_en_ctx2(MEMC6_write_mem_en_ctx2),
.mem_en_ctx2(MEMC6_mem_en_ctx2));

defparam MEMC6.DATA_WIDTH = 32;
defparam MEMC6.ADDR_WIDTH = 6;
defparam MEMC6.STRIDE_WIDTH = 1;
wire MEMC7_valid_ctx1;
wire MEMC7_valid_ctx2;
wire [31:0] MEMC7_data_from_Core;
wire [31:0] MEMC7_data_to_Core;
wire [5:0] MEMC7_addr_out_ctx1;
wire MEMC7_write_en_ctx1;
wire MEMC7_write_mem_en_ctx1;
wire MEMC7_mem_en_ctx1;
wire [5:0] MEMC7_start_addr_ctx1;
wire [0:0] MEMC7_stride_ctx1;
wire [5:0] MEMC7_addr_out_ctx2;
wire MEMC7_write_en_ctx2;
wire MEMC7_write_mem_en_ctx2;
wire MEMC7_mem_en_ctx2;
wire [5:0] MEMC7_start_addr_ctx2;
wire [0:0] MEMC7_stride_ctx2;
wire [31:0] MEMC7_data_in_ctx1;
wire [31:0] MEMC7_data_in_ctx2;
wire [31:0] MEMC7_data_out_ctx1;
wire [31:0] MEMC7_data_out_ctx2;
wire [63:0] MEMC7_burst_count_ctx1;
wire [63:0] MEMC7_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC7(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC7_data_from_Core),
.data_to_Core(MEMC7_data_to_Core),
.valid_ctx1(MEMC7_valid_ctx1),
.addr_out_ctx1(MEMC7_addr_out_ctx1),
.write_en_ctx1(MEMC7_write_en_ctx1),
.start_addr_ctx1(MEMC7_start_addr_ctx1),
.stride_ctx1(MEMC7_stride_ctx1),
.burst_count_ctx1(MEMC7_burst_count_ctx1),
.valid_ctx2(MEMC7_valid_ctx2),
.addr_out_ctx2(MEMC7_addr_out_ctx2),
.write_en_ctx2(MEMC7_write_en_ctx2),
.start_addr_ctx2(MEMC7_start_addr_ctx2),
.stride_ctx2(MEMC7_stride_ctx2),
.burst_count_ctx2(MEMC7_burst_count_ctx2),
.data_in_ctx1(MEMC7_data_in_ctx1),
.data_in_ctx2(MEMC7_data_in_ctx2),
.data_out_ctx1(MEMC7_data_out_ctx1),
.data_out_ctx2(MEMC7_data_out_ctx2),
.write_mem_en_ctx1(MEMC7_write_mem_en_ctx1),
.mem_en_ctx1(MEMC7_mem_en_ctx1),.write_mem_en_ctx2(MEMC7_write_mem_en_ctx2),
.mem_en_ctx2(MEMC7_mem_en_ctx2));

defparam MEMC7.DATA_WIDTH = 32;
defparam MEMC7.ADDR_WIDTH = 6;
defparam MEMC7.STRIDE_WIDTH = 1;
wire MEMC8_valid_ctx1;
wire MEMC8_valid_ctx2;
wire [31:0] MEMC8_data_from_Core;
wire [31:0] MEMC8_data_to_Core;
wire [5:0] MEMC8_addr_out_ctx1;
wire MEMC8_write_en_ctx1;
wire MEMC8_write_mem_en_ctx1;
wire MEMC8_mem_en_ctx1;
wire [5:0] MEMC8_start_addr_ctx1;
wire [0:0] MEMC8_stride_ctx1;
wire [5:0] MEMC8_addr_out_ctx2;
wire MEMC8_write_en_ctx2;
wire MEMC8_write_mem_en_ctx2;
wire MEMC8_mem_en_ctx2;
wire [5:0] MEMC8_start_addr_ctx2;
wire [0:0] MEMC8_stride_ctx2;
wire [31:0] MEMC8_data_in_ctx1;
wire [31:0] MEMC8_data_in_ctx2;
wire [31:0] MEMC8_data_out_ctx1;
wire [31:0] MEMC8_data_out_ctx2;
wire [63:0] MEMC8_burst_count_ctx1;
wire [63:0] MEMC8_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC8(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC8_data_from_Core),
.data_to_Core(MEMC8_data_to_Core),
.valid_ctx1(MEMC8_valid_ctx1),
.addr_out_ctx1(MEMC8_addr_out_ctx1),
.write_en_ctx1(MEMC8_write_en_ctx1),
.start_addr_ctx1(MEMC8_start_addr_ctx1),
.stride_ctx1(MEMC8_stride_ctx1),
.burst_count_ctx1(MEMC8_burst_count_ctx1),
.valid_ctx2(MEMC8_valid_ctx2),
.addr_out_ctx2(MEMC8_addr_out_ctx2),
.write_en_ctx2(MEMC8_write_en_ctx2),
.start_addr_ctx2(MEMC8_start_addr_ctx2),
.stride_ctx2(MEMC8_stride_ctx2),
.burst_count_ctx2(MEMC8_burst_count_ctx2),
.data_in_ctx1(MEMC8_data_in_ctx1),
.data_in_ctx2(MEMC8_data_in_ctx2),
.data_out_ctx1(MEMC8_data_out_ctx1),
.data_out_ctx2(MEMC8_data_out_ctx2),
.write_mem_en_ctx1(MEMC8_write_mem_en_ctx1),
.mem_en_ctx1(MEMC8_mem_en_ctx1),.write_mem_en_ctx2(MEMC8_write_mem_en_ctx2),
.mem_en_ctx2(MEMC8_mem_en_ctx2));

defparam MEMC8.DATA_WIDTH = 32;
defparam MEMC8.ADDR_WIDTH = 6;
defparam MEMC8.STRIDE_WIDTH = 1;
wire MEMC9_valid_ctx1;
wire MEMC9_valid_ctx2;
wire [31:0] MEMC9_data_from_Core;
wire [31:0] MEMC9_data_to_Core;
wire [5:0] MEMC9_addr_out_ctx1;
wire MEMC9_write_en_ctx1;
wire MEMC9_write_mem_en_ctx1;
wire MEMC9_mem_en_ctx1;
wire [5:0] MEMC9_start_addr_ctx1;
wire [0:0] MEMC9_stride_ctx1;
wire [5:0] MEMC9_addr_out_ctx2;
wire MEMC9_write_en_ctx2;
wire MEMC9_write_mem_en_ctx2;
wire MEMC9_mem_en_ctx2;
wire [5:0] MEMC9_start_addr_ctx2;
wire [0:0] MEMC9_stride_ctx2;
wire [31:0] MEMC9_data_in_ctx1;
wire [31:0] MEMC9_data_in_ctx2;
wire [31:0] MEMC9_data_out_ctx1;
wire [31:0] MEMC9_data_out_ctx2;
wire [63:0] MEMC9_burst_count_ctx1;
wire [63:0] MEMC9_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC9(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC9_data_from_Core),
.data_to_Core(MEMC9_data_to_Core),
.valid_ctx1(MEMC9_valid_ctx1),
.addr_out_ctx1(MEMC9_addr_out_ctx1),
.write_en_ctx1(MEMC9_write_en_ctx1),
.start_addr_ctx1(MEMC9_start_addr_ctx1),
.stride_ctx1(MEMC9_stride_ctx1),
.burst_count_ctx1(MEMC9_burst_count_ctx1),
.valid_ctx2(MEMC9_valid_ctx2),
.addr_out_ctx2(MEMC9_addr_out_ctx2),
.write_en_ctx2(MEMC9_write_en_ctx2),
.start_addr_ctx2(MEMC9_start_addr_ctx2),
.stride_ctx2(MEMC9_stride_ctx2),
.burst_count_ctx2(MEMC9_burst_count_ctx2),
.data_in_ctx1(MEMC9_data_in_ctx1),
.data_in_ctx2(MEMC9_data_in_ctx2),
.data_out_ctx1(MEMC9_data_out_ctx1),
.data_out_ctx2(MEMC9_data_out_ctx2),
.write_mem_en_ctx1(MEMC9_write_mem_en_ctx1),
.mem_en_ctx1(MEMC9_mem_en_ctx1),.write_mem_en_ctx2(MEMC9_write_mem_en_ctx2),
.mem_en_ctx2(MEMC9_mem_en_ctx2));

defparam MEMC9.DATA_WIDTH = 32;
defparam MEMC9.ADDR_WIDTH = 6;
defparam MEMC9.STRIDE_WIDTH = 1;
wire MEMC10_valid_ctx1;
wire MEMC10_valid_ctx2;
wire [31:0] MEMC10_data_from_Core;
wire [31:0] MEMC10_data_to_Core;
wire [5:0] MEMC10_addr_out_ctx1;
wire MEMC10_write_en_ctx1;
wire MEMC10_write_mem_en_ctx1;
wire MEMC10_mem_en_ctx1;
wire [5:0] MEMC10_start_addr_ctx1;
wire [0:0] MEMC10_stride_ctx1;
wire [5:0] MEMC10_addr_out_ctx2;
wire MEMC10_write_en_ctx2;
wire MEMC10_write_mem_en_ctx2;
wire MEMC10_mem_en_ctx2;
wire [5:0] MEMC10_start_addr_ctx2;
wire [0:0] MEMC10_stride_ctx2;
wire [31:0] MEMC10_data_in_ctx1;
wire [31:0] MEMC10_data_in_ctx2;
wire [31:0] MEMC10_data_out_ctx1;
wire [31:0] MEMC10_data_out_ctx2;
wire [63:0] MEMC10_burst_count_ctx1;
wire [63:0] MEMC10_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC10(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC10_data_from_Core),
.data_to_Core(MEMC10_data_to_Core),
.valid_ctx1(MEMC10_valid_ctx1),
.addr_out_ctx1(MEMC10_addr_out_ctx1),
.write_en_ctx1(MEMC10_write_en_ctx1),
.start_addr_ctx1(MEMC10_start_addr_ctx1),
.stride_ctx1(MEMC10_stride_ctx1),
.burst_count_ctx1(MEMC10_burst_count_ctx1),
.valid_ctx2(MEMC10_valid_ctx2),
.addr_out_ctx2(MEMC10_addr_out_ctx2),
.write_en_ctx2(MEMC10_write_en_ctx2),
.start_addr_ctx2(MEMC10_start_addr_ctx2),
.stride_ctx2(MEMC10_stride_ctx2),
.burst_count_ctx2(MEMC10_burst_count_ctx2),
.data_in_ctx1(MEMC10_data_in_ctx1),
.data_in_ctx2(MEMC10_data_in_ctx2),
.data_out_ctx1(MEMC10_data_out_ctx1),
.data_out_ctx2(MEMC10_data_out_ctx2),
.write_mem_en_ctx1(MEMC10_write_mem_en_ctx1),
.mem_en_ctx1(MEMC10_mem_en_ctx1),.write_mem_en_ctx2(MEMC10_write_mem_en_ctx2),
.mem_en_ctx2(MEMC10_mem_en_ctx2));

defparam MEMC10.DATA_WIDTH = 32;
defparam MEMC10.ADDR_WIDTH = 6;
defparam MEMC10.STRIDE_WIDTH = 1;
wire MEMC11_valid_ctx1;
wire MEMC11_valid_ctx2;
wire [31:0] MEMC11_data_from_Core;
wire [31:0] MEMC11_data_to_Core;
wire [5:0] MEMC11_addr_out_ctx1;
wire MEMC11_write_en_ctx1;
wire MEMC11_write_mem_en_ctx1;
wire MEMC11_mem_en_ctx1;
wire [5:0] MEMC11_start_addr_ctx1;
wire [0:0] MEMC11_stride_ctx1;
wire [5:0] MEMC11_addr_out_ctx2;
wire MEMC11_write_en_ctx2;
wire MEMC11_write_mem_en_ctx2;
wire MEMC11_mem_en_ctx2;
wire [5:0] MEMC11_start_addr_ctx2;
wire [0:0] MEMC11_stride_ctx2;
wire [31:0] MEMC11_data_in_ctx1;
wire [31:0] MEMC11_data_in_ctx2;
wire [31:0] MEMC11_data_out_ctx1;
wire [31:0] MEMC11_data_out_ctx2;
wire [63:0] MEMC11_burst_count_ctx1;
wire [63:0] MEMC11_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC11(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC11_data_from_Core),
.data_to_Core(MEMC11_data_to_Core),
.valid_ctx1(MEMC11_valid_ctx1),
.addr_out_ctx1(MEMC11_addr_out_ctx1),
.write_en_ctx1(MEMC11_write_en_ctx1),
.start_addr_ctx1(MEMC11_start_addr_ctx1),
.stride_ctx1(MEMC11_stride_ctx1),
.burst_count_ctx1(MEMC11_burst_count_ctx1),
.valid_ctx2(MEMC11_valid_ctx2),
.addr_out_ctx2(MEMC11_addr_out_ctx2),
.write_en_ctx2(MEMC11_write_en_ctx2),
.start_addr_ctx2(MEMC11_start_addr_ctx2),
.stride_ctx2(MEMC11_stride_ctx2),
.burst_count_ctx2(MEMC11_burst_count_ctx2),
.data_in_ctx1(MEMC11_data_in_ctx1),
.data_in_ctx2(MEMC11_data_in_ctx2),
.data_out_ctx1(MEMC11_data_out_ctx1),
.data_out_ctx2(MEMC11_data_out_ctx2),
.write_mem_en_ctx1(MEMC11_write_mem_en_ctx1),
.mem_en_ctx1(MEMC11_mem_en_ctx1),.write_mem_en_ctx2(MEMC11_write_mem_en_ctx2),
.mem_en_ctx2(MEMC11_mem_en_ctx2));

defparam MEMC11.DATA_WIDTH = 32;
defparam MEMC11.ADDR_WIDTH = 6;
defparam MEMC11.STRIDE_WIDTH = 1;
wire MEMC12_valid_ctx1;
wire MEMC12_valid_ctx2;
wire [31:0] MEMC12_data_from_Core;
wire [31:0] MEMC12_data_to_Core;
wire [5:0] MEMC12_addr_out_ctx1;
wire MEMC12_write_en_ctx1;
wire MEMC12_write_mem_en_ctx1;
wire MEMC12_mem_en_ctx1;
wire [5:0] MEMC12_start_addr_ctx1;
wire [0:0] MEMC12_stride_ctx1;
wire [5:0] MEMC12_addr_out_ctx2;
wire MEMC12_write_en_ctx2;
wire MEMC12_write_mem_en_ctx2;
wire MEMC12_mem_en_ctx2;
wire [5:0] MEMC12_start_addr_ctx2;
wire [0:0] MEMC12_stride_ctx2;
wire [31:0] MEMC12_data_in_ctx1;
wire [31:0] MEMC12_data_in_ctx2;
wire [31:0] MEMC12_data_out_ctx1;
wire [31:0] MEMC12_data_out_ctx2;
wire [63:0] MEMC12_burst_count_ctx1;
wire [63:0] MEMC12_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC12(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC12_data_from_Core),
.data_to_Core(MEMC12_data_to_Core),
.valid_ctx1(MEMC12_valid_ctx1),
.addr_out_ctx1(MEMC12_addr_out_ctx1),
.write_en_ctx1(MEMC12_write_en_ctx1),
.start_addr_ctx1(MEMC12_start_addr_ctx1),
.stride_ctx1(MEMC12_stride_ctx1),
.burst_count_ctx1(MEMC12_burst_count_ctx1),
.valid_ctx2(MEMC12_valid_ctx2),
.addr_out_ctx2(MEMC12_addr_out_ctx2),
.write_en_ctx2(MEMC12_write_en_ctx2),
.start_addr_ctx2(MEMC12_start_addr_ctx2),
.stride_ctx2(MEMC12_stride_ctx2),
.burst_count_ctx2(MEMC12_burst_count_ctx2),
.data_in_ctx1(MEMC12_data_in_ctx1),
.data_in_ctx2(MEMC12_data_in_ctx2),
.data_out_ctx1(MEMC12_data_out_ctx1),
.data_out_ctx2(MEMC12_data_out_ctx2),
.write_mem_en_ctx1(MEMC12_write_mem_en_ctx1),
.mem_en_ctx1(MEMC12_mem_en_ctx1),.write_mem_en_ctx2(MEMC12_write_mem_en_ctx2),
.mem_en_ctx2(MEMC12_mem_en_ctx2));

defparam MEMC12.DATA_WIDTH = 32;
defparam MEMC12.ADDR_WIDTH = 6;
defparam MEMC12.STRIDE_WIDTH = 1;
wire MEMC13_valid_ctx1;
wire MEMC13_valid_ctx2;
wire [31:0] MEMC13_data_from_Core;
wire [31:0] MEMC13_data_to_Core;
wire [5:0] MEMC13_addr_out_ctx1;
wire MEMC13_write_en_ctx1;
wire MEMC13_write_mem_en_ctx1;
wire MEMC13_mem_en_ctx1;
wire [5:0] MEMC13_start_addr_ctx1;
wire [0:0] MEMC13_stride_ctx1;
wire [5:0] MEMC13_addr_out_ctx2;
wire MEMC13_write_en_ctx2;
wire MEMC13_write_mem_en_ctx2;
wire MEMC13_mem_en_ctx2;
wire [5:0] MEMC13_start_addr_ctx2;
wire [0:0] MEMC13_stride_ctx2;
wire [31:0] MEMC13_data_in_ctx1;
wire [31:0] MEMC13_data_in_ctx2;
wire [31:0] MEMC13_data_out_ctx1;
wire [31:0] MEMC13_data_out_ctx2;
wire [63:0] MEMC13_burst_count_ctx1;
wire [63:0] MEMC13_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC13(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC13_data_from_Core),
.data_to_Core(MEMC13_data_to_Core),
.valid_ctx1(MEMC13_valid_ctx1),
.addr_out_ctx1(MEMC13_addr_out_ctx1),
.write_en_ctx1(MEMC13_write_en_ctx1),
.start_addr_ctx1(MEMC13_start_addr_ctx1),
.stride_ctx1(MEMC13_stride_ctx1),
.burst_count_ctx1(MEMC13_burst_count_ctx1),
.valid_ctx2(MEMC13_valid_ctx2),
.addr_out_ctx2(MEMC13_addr_out_ctx2),
.write_en_ctx2(MEMC13_write_en_ctx2),
.start_addr_ctx2(MEMC13_start_addr_ctx2),
.stride_ctx2(MEMC13_stride_ctx2),
.burst_count_ctx2(MEMC13_burst_count_ctx2),
.data_in_ctx1(MEMC13_data_in_ctx1),
.data_in_ctx2(MEMC13_data_in_ctx2),
.data_out_ctx1(MEMC13_data_out_ctx1),
.data_out_ctx2(MEMC13_data_out_ctx2),
.write_mem_en_ctx1(MEMC13_write_mem_en_ctx1),
.mem_en_ctx1(MEMC13_mem_en_ctx1),.write_mem_en_ctx2(MEMC13_write_mem_en_ctx2),
.mem_en_ctx2(MEMC13_mem_en_ctx2));

defparam MEMC13.DATA_WIDTH = 32;
defparam MEMC13.ADDR_WIDTH = 6;
defparam MEMC13.STRIDE_WIDTH = 1;
wire MEMC14_valid_ctx1;
wire MEMC14_valid_ctx2;
wire [31:0] MEMC14_data_from_Core;
wire [31:0] MEMC14_data_to_Core;
wire [5:0] MEMC14_addr_out_ctx1;
wire MEMC14_write_en_ctx1;
wire MEMC14_write_mem_en_ctx1;
wire MEMC14_mem_en_ctx1;
wire [5:0] MEMC14_start_addr_ctx1;
wire [0:0] MEMC14_stride_ctx1;
wire [5:0] MEMC14_addr_out_ctx2;
wire MEMC14_write_en_ctx2;
wire MEMC14_write_mem_en_ctx2;
wire MEMC14_mem_en_ctx2;
wire [5:0] MEMC14_start_addr_ctx2;
wire [0:0] MEMC14_stride_ctx2;
wire [31:0] MEMC14_data_in_ctx1;
wire [31:0] MEMC14_data_in_ctx2;
wire [31:0] MEMC14_data_out_ctx1;
wire [31:0] MEMC14_data_out_ctx2;
wire [63:0] MEMC14_burst_count_ctx1;
wire [63:0] MEMC14_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC14(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC14_data_from_Core),
.data_to_Core(MEMC14_data_to_Core),
.valid_ctx1(MEMC14_valid_ctx1),
.addr_out_ctx1(MEMC14_addr_out_ctx1),
.write_en_ctx1(MEMC14_write_en_ctx1),
.start_addr_ctx1(MEMC14_start_addr_ctx1),
.stride_ctx1(MEMC14_stride_ctx1),
.burst_count_ctx1(MEMC14_burst_count_ctx1),
.valid_ctx2(MEMC14_valid_ctx2),
.addr_out_ctx2(MEMC14_addr_out_ctx2),
.write_en_ctx2(MEMC14_write_en_ctx2),
.start_addr_ctx2(MEMC14_start_addr_ctx2),
.stride_ctx2(MEMC14_stride_ctx2),
.burst_count_ctx2(MEMC14_burst_count_ctx2),
.data_in_ctx1(MEMC14_data_in_ctx1),
.data_in_ctx2(MEMC14_data_in_ctx2),
.data_out_ctx1(MEMC14_data_out_ctx1),
.data_out_ctx2(MEMC14_data_out_ctx2),
.write_mem_en_ctx1(MEMC14_write_mem_en_ctx1),
.mem_en_ctx1(MEMC14_mem_en_ctx1),.write_mem_en_ctx2(MEMC14_write_mem_en_ctx2),
.mem_en_ctx2(MEMC14_mem_en_ctx2));

defparam MEMC14.DATA_WIDTH = 32;
defparam MEMC14.ADDR_WIDTH = 6;
defparam MEMC14.STRIDE_WIDTH = 1;
wire MEMC15_valid_ctx1;
wire MEMC15_valid_ctx2;
wire [31:0] MEMC15_data_from_Core;
wire [31:0] MEMC15_data_to_Core;
wire [5:0] MEMC15_addr_out_ctx1;
wire MEMC15_write_en_ctx1;
wire MEMC15_write_mem_en_ctx1;
wire MEMC15_mem_en_ctx1;
wire [5:0] MEMC15_start_addr_ctx1;
wire [0:0] MEMC15_stride_ctx1;
wire [5:0] MEMC15_addr_out_ctx2;
wire MEMC15_write_en_ctx2;
wire MEMC15_write_mem_en_ctx2;
wire MEMC15_mem_en_ctx2;
wire [5:0] MEMC15_start_addr_ctx2;
wire [0:0] MEMC15_stride_ctx2;
wire [31:0] MEMC15_data_in_ctx1;
wire [31:0] MEMC15_data_in_ctx2;
wire [31:0] MEMC15_data_out_ctx1;
wire [31:0] MEMC15_data_out_ctx2;
wire [63:0] MEMC15_burst_count_ctx1;
wire [63:0] MEMC15_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC15(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC15_data_from_Core),
.data_to_Core(MEMC15_data_to_Core),
.valid_ctx1(MEMC15_valid_ctx1),
.addr_out_ctx1(MEMC15_addr_out_ctx1),
.write_en_ctx1(MEMC15_write_en_ctx1),
.start_addr_ctx1(MEMC15_start_addr_ctx1),
.stride_ctx1(MEMC15_stride_ctx1),
.burst_count_ctx1(MEMC15_burst_count_ctx1),
.valid_ctx2(MEMC15_valid_ctx2),
.addr_out_ctx2(MEMC15_addr_out_ctx2),
.write_en_ctx2(MEMC15_write_en_ctx2),
.start_addr_ctx2(MEMC15_start_addr_ctx2),
.stride_ctx2(MEMC15_stride_ctx2),
.burst_count_ctx2(MEMC15_burst_count_ctx2),
.data_in_ctx1(MEMC15_data_in_ctx1),
.data_in_ctx2(MEMC15_data_in_ctx2),
.data_out_ctx1(MEMC15_data_out_ctx1),
.data_out_ctx2(MEMC15_data_out_ctx2),
.write_mem_en_ctx1(MEMC15_write_mem_en_ctx1),
.mem_en_ctx1(MEMC15_mem_en_ctx1),.write_mem_en_ctx2(MEMC15_write_mem_en_ctx2),
.mem_en_ctx2(MEMC15_mem_en_ctx2));

defparam MEMC15.DATA_WIDTH = 32;
defparam MEMC15.ADDR_WIDTH = 6;
defparam MEMC15.STRIDE_WIDTH = 1;
wire MEMC16_valid_ctx1;
wire MEMC16_valid_ctx2;
wire [31:0] MEMC16_data_from_Core;
wire [31:0] MEMC16_data_to_Core;
wire [5:0] MEMC16_addr_out_ctx1;
wire MEMC16_write_en_ctx1;
wire MEMC16_write_mem_en_ctx1;
wire MEMC16_mem_en_ctx1;
wire [5:0] MEMC16_start_addr_ctx1;
wire [0:0] MEMC16_stride_ctx1;
wire [5:0] MEMC16_addr_out_ctx2;
wire MEMC16_write_en_ctx2;
wire MEMC16_write_mem_en_ctx2;
wire MEMC16_mem_en_ctx2;
wire [5:0] MEMC16_start_addr_ctx2;
wire [0:0] MEMC16_stride_ctx2;
wire [31:0] MEMC16_data_in_ctx1;
wire [31:0] MEMC16_data_in_ctx2;
wire [31:0] MEMC16_data_out_ctx1;
wire [31:0] MEMC16_data_out_ctx2;
wire [63:0] MEMC16_burst_count_ctx1;
wire [63:0] MEMC16_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC16(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC16_data_from_Core),
.data_to_Core(MEMC16_data_to_Core),
.valid_ctx1(MEMC16_valid_ctx1),
.addr_out_ctx1(MEMC16_addr_out_ctx1),
.write_en_ctx1(MEMC16_write_en_ctx1),
.start_addr_ctx1(MEMC16_start_addr_ctx1),
.stride_ctx1(MEMC16_stride_ctx1),
.burst_count_ctx1(MEMC16_burst_count_ctx1),
.valid_ctx2(MEMC16_valid_ctx2),
.addr_out_ctx2(MEMC16_addr_out_ctx2),
.write_en_ctx2(MEMC16_write_en_ctx2),
.start_addr_ctx2(MEMC16_start_addr_ctx2),
.stride_ctx2(MEMC16_stride_ctx2),
.burst_count_ctx2(MEMC16_burst_count_ctx2),
.data_in_ctx1(MEMC16_data_in_ctx1),
.data_in_ctx2(MEMC16_data_in_ctx2),
.data_out_ctx1(MEMC16_data_out_ctx1),
.data_out_ctx2(MEMC16_data_out_ctx2),
.write_mem_en_ctx1(MEMC16_write_mem_en_ctx1),
.mem_en_ctx1(MEMC16_mem_en_ctx1),.write_mem_en_ctx2(MEMC16_write_mem_en_ctx2),
.mem_en_ctx2(MEMC16_mem_en_ctx2));

defparam MEMC16.DATA_WIDTH = 32;
defparam MEMC16.ADDR_WIDTH = 6;
defparam MEMC16.STRIDE_WIDTH = 1;
wire MEMC17_valid_ctx1;
wire MEMC17_valid_ctx2;
wire [31:0] MEMC17_data_from_Core;
wire [31:0] MEMC17_data_to_Core;
wire [5:0] MEMC17_addr_out_ctx1;
wire MEMC17_write_en_ctx1;
wire MEMC17_write_mem_en_ctx1;
wire MEMC17_mem_en_ctx1;
wire [5:0] MEMC17_start_addr_ctx1;
wire [0:0] MEMC17_stride_ctx1;
wire [5:0] MEMC17_addr_out_ctx2;
wire MEMC17_write_en_ctx2;
wire MEMC17_write_mem_en_ctx2;
wire MEMC17_mem_en_ctx2;
wire [5:0] MEMC17_start_addr_ctx2;
wire [0:0] MEMC17_stride_ctx2;
wire [31:0] MEMC17_data_in_ctx1;
wire [31:0] MEMC17_data_in_ctx2;
wire [31:0] MEMC17_data_out_ctx1;
wire [31:0] MEMC17_data_out_ctx2;
wire [63:0] MEMC17_burst_count_ctx1;
wire [63:0] MEMC17_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC17(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC17_data_from_Core),
.data_to_Core(MEMC17_data_to_Core),
.valid_ctx1(MEMC17_valid_ctx1),
.addr_out_ctx1(MEMC17_addr_out_ctx1),
.write_en_ctx1(MEMC17_write_en_ctx1),
.start_addr_ctx1(MEMC17_start_addr_ctx1),
.stride_ctx1(MEMC17_stride_ctx1),
.burst_count_ctx1(MEMC17_burst_count_ctx1),
.valid_ctx2(MEMC17_valid_ctx2),
.addr_out_ctx2(MEMC17_addr_out_ctx2),
.write_en_ctx2(MEMC17_write_en_ctx2),
.start_addr_ctx2(MEMC17_start_addr_ctx2),
.stride_ctx2(MEMC17_stride_ctx2),
.burst_count_ctx2(MEMC17_burst_count_ctx2),
.data_in_ctx1(MEMC17_data_in_ctx1),
.data_in_ctx2(MEMC17_data_in_ctx2),
.data_out_ctx1(MEMC17_data_out_ctx1),
.data_out_ctx2(MEMC17_data_out_ctx2),
.write_mem_en_ctx1(MEMC17_write_mem_en_ctx1),
.mem_en_ctx1(MEMC17_mem_en_ctx1),.write_mem_en_ctx2(MEMC17_write_mem_en_ctx2),
.mem_en_ctx2(MEMC17_mem_en_ctx2));

defparam MEMC17.DATA_WIDTH = 32;
defparam MEMC17.ADDR_WIDTH = 6;
defparam MEMC17.STRIDE_WIDTH = 1;
wire MEMC18_valid_ctx1;
wire MEMC18_valid_ctx2;
wire [31:0] MEMC18_data_from_Core;
wire [31:0] MEMC18_data_to_Core;
wire [5:0] MEMC18_addr_out_ctx1;
wire MEMC18_write_en_ctx1;
wire MEMC18_write_mem_en_ctx1;
wire MEMC18_mem_en_ctx1;
wire [5:0] MEMC18_start_addr_ctx1;
wire [0:0] MEMC18_stride_ctx1;
wire [5:0] MEMC18_addr_out_ctx2;
wire MEMC18_write_en_ctx2;
wire MEMC18_write_mem_en_ctx2;
wire MEMC18_mem_en_ctx2;
wire [5:0] MEMC18_start_addr_ctx2;
wire [0:0] MEMC18_stride_ctx2;
wire [31:0] MEMC18_data_in_ctx1;
wire [31:0] MEMC18_data_in_ctx2;
wire [31:0] MEMC18_data_out_ctx1;
wire [31:0] MEMC18_data_out_ctx2;
wire [63:0] MEMC18_burst_count_ctx1;
wire [63:0] MEMC18_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC18(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC18_data_from_Core),
.data_to_Core(MEMC18_data_to_Core),
.valid_ctx1(MEMC18_valid_ctx1),
.addr_out_ctx1(MEMC18_addr_out_ctx1),
.write_en_ctx1(MEMC18_write_en_ctx1),
.start_addr_ctx1(MEMC18_start_addr_ctx1),
.stride_ctx1(MEMC18_stride_ctx1),
.burst_count_ctx1(MEMC18_burst_count_ctx1),
.valid_ctx2(MEMC18_valid_ctx2),
.addr_out_ctx2(MEMC18_addr_out_ctx2),
.write_en_ctx2(MEMC18_write_en_ctx2),
.start_addr_ctx2(MEMC18_start_addr_ctx2),
.stride_ctx2(MEMC18_stride_ctx2),
.burst_count_ctx2(MEMC18_burst_count_ctx2),
.data_in_ctx1(MEMC18_data_in_ctx1),
.data_in_ctx2(MEMC18_data_in_ctx2),
.data_out_ctx1(MEMC18_data_out_ctx1),
.data_out_ctx2(MEMC18_data_out_ctx2),
.write_mem_en_ctx1(MEMC18_write_mem_en_ctx1),
.mem_en_ctx1(MEMC18_mem_en_ctx1),.write_mem_en_ctx2(MEMC18_write_mem_en_ctx2),
.mem_en_ctx2(MEMC18_mem_en_ctx2));

defparam MEMC18.DATA_WIDTH = 32;
defparam MEMC18.ADDR_WIDTH = 6;
defparam MEMC18.STRIDE_WIDTH = 1;
wire MEMC19_valid_ctx1;
wire MEMC19_valid_ctx2;
wire [31:0] MEMC19_data_from_Core;
wire [31:0] MEMC19_data_to_Core;
wire [5:0] MEMC19_addr_out_ctx1;
wire MEMC19_write_en_ctx1;
wire MEMC19_write_mem_en_ctx1;
wire MEMC19_mem_en_ctx1;
wire [5:0] MEMC19_start_addr_ctx1;
wire [0:0] MEMC19_stride_ctx1;
wire [5:0] MEMC19_addr_out_ctx2;
wire MEMC19_write_en_ctx2;
wire MEMC19_write_mem_en_ctx2;
wire MEMC19_mem_en_ctx2;
wire [5:0] MEMC19_start_addr_ctx2;
wire [0:0] MEMC19_stride_ctx2;
wire [31:0] MEMC19_data_in_ctx1;
wire [31:0] MEMC19_data_in_ctx2;
wire [31:0] MEMC19_data_out_ctx1;
wire [31:0] MEMC19_data_out_ctx2;
wire [63:0] MEMC19_burst_count_ctx1;
wire [63:0] MEMC19_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC19(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC19_data_from_Core),
.data_to_Core(MEMC19_data_to_Core),
.valid_ctx1(MEMC19_valid_ctx1),
.addr_out_ctx1(MEMC19_addr_out_ctx1),
.write_en_ctx1(MEMC19_write_en_ctx1),
.start_addr_ctx1(MEMC19_start_addr_ctx1),
.stride_ctx1(MEMC19_stride_ctx1),
.burst_count_ctx1(MEMC19_burst_count_ctx1),
.valid_ctx2(MEMC19_valid_ctx2),
.addr_out_ctx2(MEMC19_addr_out_ctx2),
.write_en_ctx2(MEMC19_write_en_ctx2),
.start_addr_ctx2(MEMC19_start_addr_ctx2),
.stride_ctx2(MEMC19_stride_ctx2),
.burst_count_ctx2(MEMC19_burst_count_ctx2),
.data_in_ctx1(MEMC19_data_in_ctx1),
.data_in_ctx2(MEMC19_data_in_ctx2),
.data_out_ctx1(MEMC19_data_out_ctx1),
.data_out_ctx2(MEMC19_data_out_ctx2),
.write_mem_en_ctx1(MEMC19_write_mem_en_ctx1),
.mem_en_ctx1(MEMC19_mem_en_ctx1),.write_mem_en_ctx2(MEMC19_write_mem_en_ctx2),
.mem_en_ctx2(MEMC19_mem_en_ctx2));

defparam MEMC19.DATA_WIDTH = 32;
defparam MEMC19.ADDR_WIDTH = 6;
defparam MEMC19.STRIDE_WIDTH = 1;
wire MEMC20_valid_ctx1;
wire MEMC20_valid_ctx2;
wire [31:0] MEMC20_data_from_Core;
wire [31:0] MEMC20_data_to_Core;
wire [5:0] MEMC20_addr_out_ctx1;
wire MEMC20_write_en_ctx1;
wire MEMC20_write_mem_en_ctx1;
wire MEMC20_mem_en_ctx1;
wire [5:0] MEMC20_start_addr_ctx1;
wire [0:0] MEMC20_stride_ctx1;
wire [5:0] MEMC20_addr_out_ctx2;
wire MEMC20_write_en_ctx2;
wire MEMC20_write_mem_en_ctx2;
wire MEMC20_mem_en_ctx2;
wire [5:0] MEMC20_start_addr_ctx2;
wire [0:0] MEMC20_stride_ctx2;
wire [31:0] MEMC20_data_in_ctx1;
wire [31:0] MEMC20_data_in_ctx2;
wire [31:0] MEMC20_data_out_ctx1;
wire [31:0] MEMC20_data_out_ctx2;
wire [63:0] MEMC20_burst_count_ctx1;
wire [63:0] MEMC20_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC20(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC20_data_from_Core),
.data_to_Core(MEMC20_data_to_Core),
.valid_ctx1(MEMC20_valid_ctx1),
.addr_out_ctx1(MEMC20_addr_out_ctx1),
.write_en_ctx1(MEMC20_write_en_ctx1),
.start_addr_ctx1(MEMC20_start_addr_ctx1),
.stride_ctx1(MEMC20_stride_ctx1),
.burst_count_ctx1(MEMC20_burst_count_ctx1),
.valid_ctx2(MEMC20_valid_ctx2),
.addr_out_ctx2(MEMC20_addr_out_ctx2),
.write_en_ctx2(MEMC20_write_en_ctx2),
.start_addr_ctx2(MEMC20_start_addr_ctx2),
.stride_ctx2(MEMC20_stride_ctx2),
.burst_count_ctx2(MEMC20_burst_count_ctx2),
.data_in_ctx1(MEMC20_data_in_ctx1),
.data_in_ctx2(MEMC20_data_in_ctx2),
.data_out_ctx1(MEMC20_data_out_ctx1),
.data_out_ctx2(MEMC20_data_out_ctx2),
.write_mem_en_ctx1(MEMC20_write_mem_en_ctx1),
.mem_en_ctx1(MEMC20_mem_en_ctx1),.write_mem_en_ctx2(MEMC20_write_mem_en_ctx2),
.mem_en_ctx2(MEMC20_mem_en_ctx2));

defparam MEMC20.DATA_WIDTH = 32;
defparam MEMC20.ADDR_WIDTH = 6;
defparam MEMC20.STRIDE_WIDTH = 1;
wire MEMC21_valid_ctx1;
wire MEMC21_valid_ctx2;
wire [31:0] MEMC21_data_from_Core;
wire [31:0] MEMC21_data_to_Core;
wire [5:0] MEMC21_addr_out_ctx1;
wire MEMC21_write_en_ctx1;
wire MEMC21_write_mem_en_ctx1;
wire MEMC21_mem_en_ctx1;
wire [5:0] MEMC21_start_addr_ctx1;
wire [0:0] MEMC21_stride_ctx1;
wire [5:0] MEMC21_addr_out_ctx2;
wire MEMC21_write_en_ctx2;
wire MEMC21_write_mem_en_ctx2;
wire MEMC21_mem_en_ctx2;
wire [5:0] MEMC21_start_addr_ctx2;
wire [0:0] MEMC21_stride_ctx2;
wire [31:0] MEMC21_data_in_ctx1;
wire [31:0] MEMC21_data_in_ctx2;
wire [31:0] MEMC21_data_out_ctx1;
wire [31:0] MEMC21_data_out_ctx2;
wire [63:0] MEMC21_burst_count_ctx1;
wire [63:0] MEMC21_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC21(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC21_data_from_Core),
.data_to_Core(MEMC21_data_to_Core),
.valid_ctx1(MEMC21_valid_ctx1),
.addr_out_ctx1(MEMC21_addr_out_ctx1),
.write_en_ctx1(MEMC21_write_en_ctx1),
.start_addr_ctx1(MEMC21_start_addr_ctx1),
.stride_ctx1(MEMC21_stride_ctx1),
.burst_count_ctx1(MEMC21_burst_count_ctx1),
.valid_ctx2(MEMC21_valid_ctx2),
.addr_out_ctx2(MEMC21_addr_out_ctx2),
.write_en_ctx2(MEMC21_write_en_ctx2),
.start_addr_ctx2(MEMC21_start_addr_ctx2),
.stride_ctx2(MEMC21_stride_ctx2),
.burst_count_ctx2(MEMC21_burst_count_ctx2),
.data_in_ctx1(MEMC21_data_in_ctx1),
.data_in_ctx2(MEMC21_data_in_ctx2),
.data_out_ctx1(MEMC21_data_out_ctx1),
.data_out_ctx2(MEMC21_data_out_ctx2),
.write_mem_en_ctx1(MEMC21_write_mem_en_ctx1),
.mem_en_ctx1(MEMC21_mem_en_ctx1),.write_mem_en_ctx2(MEMC21_write_mem_en_ctx2),
.mem_en_ctx2(MEMC21_mem_en_ctx2));

defparam MEMC21.DATA_WIDTH = 32;
defparam MEMC21.ADDR_WIDTH = 6;
defparam MEMC21.STRIDE_WIDTH = 1;
wire MEMC22_valid_ctx1;
wire MEMC22_valid_ctx2;
wire [31:0] MEMC22_data_from_Core;
wire [31:0] MEMC22_data_to_Core;
wire [5:0] MEMC22_addr_out_ctx1;
wire MEMC22_write_en_ctx1;
wire MEMC22_write_mem_en_ctx1;
wire MEMC22_mem_en_ctx1;
wire [5:0] MEMC22_start_addr_ctx1;
wire [0:0] MEMC22_stride_ctx1;
wire [5:0] MEMC22_addr_out_ctx2;
wire MEMC22_write_en_ctx2;
wire MEMC22_write_mem_en_ctx2;
wire MEMC22_mem_en_ctx2;
wire [5:0] MEMC22_start_addr_ctx2;
wire [0:0] MEMC22_stride_ctx2;
wire [31:0] MEMC22_data_in_ctx1;
wire [31:0] MEMC22_data_in_ctx2;
wire [31:0] MEMC22_data_out_ctx1;
wire [31:0] MEMC22_data_out_ctx2;
wire [63:0] MEMC22_burst_count_ctx1;
wire [63:0] MEMC22_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC22(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC22_data_from_Core),
.data_to_Core(MEMC22_data_to_Core),
.valid_ctx1(MEMC22_valid_ctx1),
.addr_out_ctx1(MEMC22_addr_out_ctx1),
.write_en_ctx1(MEMC22_write_en_ctx1),
.start_addr_ctx1(MEMC22_start_addr_ctx1),
.stride_ctx1(MEMC22_stride_ctx1),
.burst_count_ctx1(MEMC22_burst_count_ctx1),
.valid_ctx2(MEMC22_valid_ctx2),
.addr_out_ctx2(MEMC22_addr_out_ctx2),
.write_en_ctx2(MEMC22_write_en_ctx2),
.start_addr_ctx2(MEMC22_start_addr_ctx2),
.stride_ctx2(MEMC22_stride_ctx2),
.burst_count_ctx2(MEMC22_burst_count_ctx2),
.data_in_ctx1(MEMC22_data_in_ctx1),
.data_in_ctx2(MEMC22_data_in_ctx2),
.data_out_ctx1(MEMC22_data_out_ctx1),
.data_out_ctx2(MEMC22_data_out_ctx2),
.write_mem_en_ctx1(MEMC22_write_mem_en_ctx1),
.mem_en_ctx1(MEMC22_mem_en_ctx1),.write_mem_en_ctx2(MEMC22_write_mem_en_ctx2),
.mem_en_ctx2(MEMC22_mem_en_ctx2));

defparam MEMC22.DATA_WIDTH = 32;
defparam MEMC22.ADDR_WIDTH = 6;
defparam MEMC22.STRIDE_WIDTH = 1;
wire MEMC23_valid_ctx1;
wire MEMC23_valid_ctx2;
wire [31:0] MEMC23_data_from_Core;
wire [31:0] MEMC23_data_to_Core;
wire [5:0] MEMC23_addr_out_ctx1;
wire MEMC23_write_en_ctx1;
wire MEMC23_write_mem_en_ctx1;
wire MEMC23_mem_en_ctx1;
wire [5:0] MEMC23_start_addr_ctx1;
wire [0:0] MEMC23_stride_ctx1;
wire [5:0] MEMC23_addr_out_ctx2;
wire MEMC23_write_en_ctx2;
wire MEMC23_write_mem_en_ctx2;
wire MEMC23_mem_en_ctx2;
wire [5:0] MEMC23_start_addr_ctx2;
wire [0:0] MEMC23_stride_ctx2;
wire [31:0] MEMC23_data_in_ctx1;
wire [31:0] MEMC23_data_in_ctx2;
wire [31:0] MEMC23_data_out_ctx1;
wire [31:0] MEMC23_data_out_ctx2;
wire [63:0] MEMC23_burst_count_ctx1;
wire [63:0] MEMC23_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC23(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC23_data_from_Core),
.data_to_Core(MEMC23_data_to_Core),
.valid_ctx1(MEMC23_valid_ctx1),
.addr_out_ctx1(MEMC23_addr_out_ctx1),
.write_en_ctx1(MEMC23_write_en_ctx1),
.start_addr_ctx1(MEMC23_start_addr_ctx1),
.stride_ctx1(MEMC23_stride_ctx1),
.burst_count_ctx1(MEMC23_burst_count_ctx1),
.valid_ctx2(MEMC23_valid_ctx2),
.addr_out_ctx2(MEMC23_addr_out_ctx2),
.write_en_ctx2(MEMC23_write_en_ctx2),
.start_addr_ctx2(MEMC23_start_addr_ctx2),
.stride_ctx2(MEMC23_stride_ctx2),
.burst_count_ctx2(MEMC23_burst_count_ctx2),
.data_in_ctx1(MEMC23_data_in_ctx1),
.data_in_ctx2(MEMC23_data_in_ctx2),
.data_out_ctx1(MEMC23_data_out_ctx1),
.data_out_ctx2(MEMC23_data_out_ctx2),
.write_mem_en_ctx1(MEMC23_write_mem_en_ctx1),
.mem_en_ctx1(MEMC23_mem_en_ctx1),.write_mem_en_ctx2(MEMC23_write_mem_en_ctx2),
.mem_en_ctx2(MEMC23_mem_en_ctx2));

defparam MEMC23.DATA_WIDTH = 32;
defparam MEMC23.ADDR_WIDTH = 6;
defparam MEMC23.STRIDE_WIDTH = 1;
wire MEMC24_valid_ctx1;
wire MEMC24_valid_ctx2;
wire [31:0] MEMC24_data_from_Core;
wire [31:0] MEMC24_data_to_Core;
wire [5:0] MEMC24_addr_out_ctx1;
wire MEMC24_write_en_ctx1;
wire MEMC24_write_mem_en_ctx1;
wire MEMC24_mem_en_ctx1;
wire [5:0] MEMC24_start_addr_ctx1;
wire [0:0] MEMC24_stride_ctx1;
wire [5:0] MEMC24_addr_out_ctx2;
wire MEMC24_write_en_ctx2;
wire MEMC24_write_mem_en_ctx2;
wire MEMC24_mem_en_ctx2;
wire [5:0] MEMC24_start_addr_ctx2;
wire [0:0] MEMC24_stride_ctx2;
wire [31:0] MEMC24_data_in_ctx1;
wire [31:0] MEMC24_data_in_ctx2;
wire [31:0] MEMC24_data_out_ctx1;
wire [31:0] MEMC24_data_out_ctx2;
wire [63:0] MEMC24_burst_count_ctx1;
wire [63:0] MEMC24_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC24(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC24_data_from_Core),
.data_to_Core(MEMC24_data_to_Core),
.valid_ctx1(MEMC24_valid_ctx1),
.addr_out_ctx1(MEMC24_addr_out_ctx1),
.write_en_ctx1(MEMC24_write_en_ctx1),
.start_addr_ctx1(MEMC24_start_addr_ctx1),
.stride_ctx1(MEMC24_stride_ctx1),
.burst_count_ctx1(MEMC24_burst_count_ctx1),
.valid_ctx2(MEMC24_valid_ctx2),
.addr_out_ctx2(MEMC24_addr_out_ctx2),
.write_en_ctx2(MEMC24_write_en_ctx2),
.start_addr_ctx2(MEMC24_start_addr_ctx2),
.stride_ctx2(MEMC24_stride_ctx2),
.burst_count_ctx2(MEMC24_burst_count_ctx2),
.data_in_ctx1(MEMC24_data_in_ctx1),
.data_in_ctx2(MEMC24_data_in_ctx2),
.data_out_ctx1(MEMC24_data_out_ctx1),
.data_out_ctx2(MEMC24_data_out_ctx2),
.write_mem_en_ctx1(MEMC24_write_mem_en_ctx1),
.mem_en_ctx1(MEMC24_mem_en_ctx1),.write_mem_en_ctx2(MEMC24_write_mem_en_ctx2),
.mem_en_ctx2(MEMC24_mem_en_ctx2));

defparam MEMC24.DATA_WIDTH = 32;
defparam MEMC24.ADDR_WIDTH = 6;
defparam MEMC24.STRIDE_WIDTH = 1;
wire MEMC25_valid_ctx1;
wire MEMC25_valid_ctx2;
wire [31:0] MEMC25_data_from_Core;
wire [31:0] MEMC25_data_to_Core;
wire [5:0] MEMC25_addr_out_ctx1;
wire MEMC25_write_en_ctx1;
wire MEMC25_write_mem_en_ctx1;
wire MEMC25_mem_en_ctx1;
wire [5:0] MEMC25_start_addr_ctx1;
wire [0:0] MEMC25_stride_ctx1;
wire [5:0] MEMC25_addr_out_ctx2;
wire MEMC25_write_en_ctx2;
wire MEMC25_write_mem_en_ctx2;
wire MEMC25_mem_en_ctx2;
wire [5:0] MEMC25_start_addr_ctx2;
wire [0:0] MEMC25_stride_ctx2;
wire [31:0] MEMC25_data_in_ctx1;
wire [31:0] MEMC25_data_in_ctx2;
wire [31:0] MEMC25_data_out_ctx1;
wire [31:0] MEMC25_data_out_ctx2;
wire [63:0] MEMC25_burst_count_ctx1;
wire [63:0] MEMC25_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC25(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC25_data_from_Core),
.data_to_Core(MEMC25_data_to_Core),
.valid_ctx1(MEMC25_valid_ctx1),
.addr_out_ctx1(MEMC25_addr_out_ctx1),
.write_en_ctx1(MEMC25_write_en_ctx1),
.start_addr_ctx1(MEMC25_start_addr_ctx1),
.stride_ctx1(MEMC25_stride_ctx1),
.burst_count_ctx1(MEMC25_burst_count_ctx1),
.valid_ctx2(MEMC25_valid_ctx2),
.addr_out_ctx2(MEMC25_addr_out_ctx2),
.write_en_ctx2(MEMC25_write_en_ctx2),
.start_addr_ctx2(MEMC25_start_addr_ctx2),
.stride_ctx2(MEMC25_stride_ctx2),
.burst_count_ctx2(MEMC25_burst_count_ctx2),
.data_in_ctx1(MEMC25_data_in_ctx1),
.data_in_ctx2(MEMC25_data_in_ctx2),
.data_out_ctx1(MEMC25_data_out_ctx1),
.data_out_ctx2(MEMC25_data_out_ctx2),
.write_mem_en_ctx1(MEMC25_write_mem_en_ctx1),
.mem_en_ctx1(MEMC25_mem_en_ctx1),.write_mem_en_ctx2(MEMC25_write_mem_en_ctx2),
.mem_en_ctx2(MEMC25_mem_en_ctx2));

defparam MEMC25.DATA_WIDTH = 32;
defparam MEMC25.ADDR_WIDTH = 6;
defparam MEMC25.STRIDE_WIDTH = 1;
wire MEMC26_valid_ctx1;
wire MEMC26_valid_ctx2;
wire [31:0] MEMC26_data_from_Core;
wire [31:0] MEMC26_data_to_Core;
wire [5:0] MEMC26_addr_out_ctx1;
wire MEMC26_write_en_ctx1;
wire MEMC26_write_mem_en_ctx1;
wire MEMC26_mem_en_ctx1;
wire [5:0] MEMC26_start_addr_ctx1;
wire [0:0] MEMC26_stride_ctx1;
wire [5:0] MEMC26_addr_out_ctx2;
wire MEMC26_write_en_ctx2;
wire MEMC26_write_mem_en_ctx2;
wire MEMC26_mem_en_ctx2;
wire [5:0] MEMC26_start_addr_ctx2;
wire [0:0] MEMC26_stride_ctx2;
wire [31:0] MEMC26_data_in_ctx1;
wire [31:0] MEMC26_data_in_ctx2;
wire [31:0] MEMC26_data_out_ctx1;
wire [31:0] MEMC26_data_out_ctx2;
wire [63:0] MEMC26_burst_count_ctx1;
wire [63:0] MEMC26_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC26(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC26_data_from_Core),
.data_to_Core(MEMC26_data_to_Core),
.valid_ctx1(MEMC26_valid_ctx1),
.addr_out_ctx1(MEMC26_addr_out_ctx1),
.write_en_ctx1(MEMC26_write_en_ctx1),
.start_addr_ctx1(MEMC26_start_addr_ctx1),
.stride_ctx1(MEMC26_stride_ctx1),
.burst_count_ctx1(MEMC26_burst_count_ctx1),
.valid_ctx2(MEMC26_valid_ctx2),
.addr_out_ctx2(MEMC26_addr_out_ctx2),
.write_en_ctx2(MEMC26_write_en_ctx2),
.start_addr_ctx2(MEMC26_start_addr_ctx2),
.stride_ctx2(MEMC26_stride_ctx2),
.burst_count_ctx2(MEMC26_burst_count_ctx2),
.data_in_ctx1(MEMC26_data_in_ctx1),
.data_in_ctx2(MEMC26_data_in_ctx2),
.data_out_ctx1(MEMC26_data_out_ctx1),
.data_out_ctx2(MEMC26_data_out_ctx2),
.write_mem_en_ctx1(MEMC26_write_mem_en_ctx1),
.mem_en_ctx1(MEMC26_mem_en_ctx1),.write_mem_en_ctx2(MEMC26_write_mem_en_ctx2),
.mem_en_ctx2(MEMC26_mem_en_ctx2));

defparam MEMC26.DATA_WIDTH = 32;
defparam MEMC26.ADDR_WIDTH = 6;
defparam MEMC26.STRIDE_WIDTH = 1;
wire MEMC27_valid_ctx1;
wire MEMC27_valid_ctx2;
wire [31:0] MEMC27_data_from_Core;
wire [31:0] MEMC27_data_to_Core;
wire [5:0] MEMC27_addr_out_ctx1;
wire MEMC27_write_en_ctx1;
wire MEMC27_write_mem_en_ctx1;
wire MEMC27_mem_en_ctx1;
wire [5:0] MEMC27_start_addr_ctx1;
wire [0:0] MEMC27_stride_ctx1;
wire [5:0] MEMC27_addr_out_ctx2;
wire MEMC27_write_en_ctx2;
wire MEMC27_write_mem_en_ctx2;
wire MEMC27_mem_en_ctx2;
wire [5:0] MEMC27_start_addr_ctx2;
wire [0:0] MEMC27_stride_ctx2;
wire [31:0] MEMC27_data_in_ctx1;
wire [31:0] MEMC27_data_in_ctx2;
wire [31:0] MEMC27_data_out_ctx1;
wire [31:0] MEMC27_data_out_ctx2;
wire [63:0] MEMC27_burst_count_ctx1;
wire [63:0] MEMC27_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC27(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC27_data_from_Core),
.data_to_Core(MEMC27_data_to_Core),
.valid_ctx1(MEMC27_valid_ctx1),
.addr_out_ctx1(MEMC27_addr_out_ctx1),
.write_en_ctx1(MEMC27_write_en_ctx1),
.start_addr_ctx1(MEMC27_start_addr_ctx1),
.stride_ctx1(MEMC27_stride_ctx1),
.burst_count_ctx1(MEMC27_burst_count_ctx1),
.valid_ctx2(MEMC27_valid_ctx2),
.addr_out_ctx2(MEMC27_addr_out_ctx2),
.write_en_ctx2(MEMC27_write_en_ctx2),
.start_addr_ctx2(MEMC27_start_addr_ctx2),
.stride_ctx2(MEMC27_stride_ctx2),
.burst_count_ctx2(MEMC27_burst_count_ctx2),
.data_in_ctx1(MEMC27_data_in_ctx1),
.data_in_ctx2(MEMC27_data_in_ctx2),
.data_out_ctx1(MEMC27_data_out_ctx1),
.data_out_ctx2(MEMC27_data_out_ctx2),
.write_mem_en_ctx1(MEMC27_write_mem_en_ctx1),
.mem_en_ctx1(MEMC27_mem_en_ctx1),.write_mem_en_ctx2(MEMC27_write_mem_en_ctx2),
.mem_en_ctx2(MEMC27_mem_en_ctx2));

defparam MEMC27.DATA_WIDTH = 32;
defparam MEMC27.ADDR_WIDTH = 6;
defparam MEMC27.STRIDE_WIDTH = 1;
wire MEMC28_valid_ctx1;
wire MEMC28_valid_ctx2;
wire [31:0] MEMC28_data_from_Core;
wire [31:0] MEMC28_data_to_Core;
wire [5:0] MEMC28_addr_out_ctx1;
wire MEMC28_write_en_ctx1;
wire MEMC28_write_mem_en_ctx1;
wire MEMC28_mem_en_ctx1;
wire [5:0] MEMC28_start_addr_ctx1;
wire [0:0] MEMC28_stride_ctx1;
wire [5:0] MEMC28_addr_out_ctx2;
wire MEMC28_write_en_ctx2;
wire MEMC28_write_mem_en_ctx2;
wire MEMC28_mem_en_ctx2;
wire [5:0] MEMC28_start_addr_ctx2;
wire [0:0] MEMC28_stride_ctx2;
wire [31:0] MEMC28_data_in_ctx1;
wire [31:0] MEMC28_data_in_ctx2;
wire [31:0] MEMC28_data_out_ctx1;
wire [31:0] MEMC28_data_out_ctx2;
wire [63:0] MEMC28_burst_count_ctx1;
wire [63:0] MEMC28_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC28(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC28_data_from_Core),
.data_to_Core(MEMC28_data_to_Core),
.valid_ctx1(MEMC28_valid_ctx1),
.addr_out_ctx1(MEMC28_addr_out_ctx1),
.write_en_ctx1(MEMC28_write_en_ctx1),
.start_addr_ctx1(MEMC28_start_addr_ctx1),
.stride_ctx1(MEMC28_stride_ctx1),
.burst_count_ctx1(MEMC28_burst_count_ctx1),
.valid_ctx2(MEMC28_valid_ctx2),
.addr_out_ctx2(MEMC28_addr_out_ctx2),
.write_en_ctx2(MEMC28_write_en_ctx2),
.start_addr_ctx2(MEMC28_start_addr_ctx2),
.stride_ctx2(MEMC28_stride_ctx2),
.burst_count_ctx2(MEMC28_burst_count_ctx2),
.data_in_ctx1(MEMC28_data_in_ctx1),
.data_in_ctx2(MEMC28_data_in_ctx2),
.data_out_ctx1(MEMC28_data_out_ctx1),
.data_out_ctx2(MEMC28_data_out_ctx2),
.write_mem_en_ctx1(MEMC28_write_mem_en_ctx1),
.mem_en_ctx1(MEMC28_mem_en_ctx1),.write_mem_en_ctx2(MEMC28_write_mem_en_ctx2),
.mem_en_ctx2(MEMC28_mem_en_ctx2));

defparam MEMC28.DATA_WIDTH = 32;
defparam MEMC28.ADDR_WIDTH = 6;
defparam MEMC28.STRIDE_WIDTH = 1;
wire MEMC29_valid_ctx1;
wire MEMC29_valid_ctx2;
wire [31:0] MEMC29_data_from_Core;
wire [31:0] MEMC29_data_to_Core;
wire [5:0] MEMC29_addr_out_ctx1;
wire MEMC29_write_en_ctx1;
wire MEMC29_write_mem_en_ctx1;
wire MEMC29_mem_en_ctx1;
wire [5:0] MEMC29_start_addr_ctx1;
wire [0:0] MEMC29_stride_ctx1;
wire [5:0] MEMC29_addr_out_ctx2;
wire MEMC29_write_en_ctx2;
wire MEMC29_write_mem_en_ctx2;
wire MEMC29_mem_en_ctx2;
wire [5:0] MEMC29_start_addr_ctx2;
wire [0:0] MEMC29_stride_ctx2;
wire [31:0] MEMC29_data_in_ctx1;
wire [31:0] MEMC29_data_in_ctx2;
wire [31:0] MEMC29_data_out_ctx1;
wire [31:0] MEMC29_data_out_ctx2;
wire [63:0] MEMC29_burst_count_ctx1;
wire [63:0] MEMC29_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC29(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC29_data_from_Core),
.data_to_Core(MEMC29_data_to_Core),
.valid_ctx1(MEMC29_valid_ctx1),
.addr_out_ctx1(MEMC29_addr_out_ctx1),
.write_en_ctx1(MEMC29_write_en_ctx1),
.start_addr_ctx1(MEMC29_start_addr_ctx1),
.stride_ctx1(MEMC29_stride_ctx1),
.burst_count_ctx1(MEMC29_burst_count_ctx1),
.valid_ctx2(MEMC29_valid_ctx2),
.addr_out_ctx2(MEMC29_addr_out_ctx2),
.write_en_ctx2(MEMC29_write_en_ctx2),
.start_addr_ctx2(MEMC29_start_addr_ctx2),
.stride_ctx2(MEMC29_stride_ctx2),
.burst_count_ctx2(MEMC29_burst_count_ctx2),
.data_in_ctx1(MEMC29_data_in_ctx1),
.data_in_ctx2(MEMC29_data_in_ctx2),
.data_out_ctx1(MEMC29_data_out_ctx1),
.data_out_ctx2(MEMC29_data_out_ctx2),
.write_mem_en_ctx1(MEMC29_write_mem_en_ctx1),
.mem_en_ctx1(MEMC29_mem_en_ctx1),.write_mem_en_ctx2(MEMC29_write_mem_en_ctx2),
.mem_en_ctx2(MEMC29_mem_en_ctx2));

defparam MEMC29.DATA_WIDTH = 32;
defparam MEMC29.ADDR_WIDTH = 6;
defparam MEMC29.STRIDE_WIDTH = 1;
wire MEMC30_valid_ctx1;
wire MEMC30_valid_ctx2;
wire [31:0] MEMC30_data_from_Core;
wire [31:0] MEMC30_data_to_Core;
wire [5:0] MEMC30_addr_out_ctx1;
wire MEMC30_write_en_ctx1;
wire MEMC30_write_mem_en_ctx1;
wire MEMC30_mem_en_ctx1;
wire [5:0] MEMC30_start_addr_ctx1;
wire [0:0] MEMC30_stride_ctx1;
wire [5:0] MEMC30_addr_out_ctx2;
wire MEMC30_write_en_ctx2;
wire MEMC30_write_mem_en_ctx2;
wire MEMC30_mem_en_ctx2;
wire [5:0] MEMC30_start_addr_ctx2;
wire [0:0] MEMC30_stride_ctx2;
wire [31:0] MEMC30_data_in_ctx1;
wire [31:0] MEMC30_data_in_ctx2;
wire [31:0] MEMC30_data_out_ctx1;
wire [31:0] MEMC30_data_out_ctx2;
wire [63:0] MEMC30_burst_count_ctx1;
wire [63:0] MEMC30_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC30(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC30_data_from_Core),
.data_to_Core(MEMC30_data_to_Core),
.valid_ctx1(MEMC30_valid_ctx1),
.addr_out_ctx1(MEMC30_addr_out_ctx1),
.write_en_ctx1(MEMC30_write_en_ctx1),
.start_addr_ctx1(MEMC30_start_addr_ctx1),
.stride_ctx1(MEMC30_stride_ctx1),
.burst_count_ctx1(MEMC30_burst_count_ctx1),
.valid_ctx2(MEMC30_valid_ctx2),
.addr_out_ctx2(MEMC30_addr_out_ctx2),
.write_en_ctx2(MEMC30_write_en_ctx2),
.start_addr_ctx2(MEMC30_start_addr_ctx2),
.stride_ctx2(MEMC30_stride_ctx2),
.burst_count_ctx2(MEMC30_burst_count_ctx2),
.data_in_ctx1(MEMC30_data_in_ctx1),
.data_in_ctx2(MEMC30_data_in_ctx2),
.data_out_ctx1(MEMC30_data_out_ctx1),
.data_out_ctx2(MEMC30_data_out_ctx2),
.write_mem_en_ctx1(MEMC30_write_mem_en_ctx1),
.mem_en_ctx1(MEMC30_mem_en_ctx1),.write_mem_en_ctx2(MEMC30_write_mem_en_ctx2),
.mem_en_ctx2(MEMC30_mem_en_ctx2));

defparam MEMC30.DATA_WIDTH = 32;
defparam MEMC30.ADDR_WIDTH = 6;
defparam MEMC30.STRIDE_WIDTH = 1;
wire MEMC31_valid_ctx1;
wire MEMC31_valid_ctx2;
wire [31:0] MEMC31_data_from_Core;
wire [31:0] MEMC31_data_to_Core;
wire [5:0] MEMC31_addr_out_ctx1;
wire MEMC31_write_en_ctx1;
wire MEMC31_write_mem_en_ctx1;
wire MEMC31_mem_en_ctx1;
wire [5:0] MEMC31_start_addr_ctx1;
wire [0:0] MEMC31_stride_ctx1;
wire [5:0] MEMC31_addr_out_ctx2;
wire MEMC31_write_en_ctx2;
wire MEMC31_write_mem_en_ctx2;
wire MEMC31_mem_en_ctx2;
wire [5:0] MEMC31_start_addr_ctx2;
wire [0:0] MEMC31_stride_ctx2;
wire [31:0] MEMC31_data_in_ctx1;
wire [31:0] MEMC31_data_in_ctx2;
wire [31:0] MEMC31_data_out_ctx1;
wire [31:0] MEMC31_data_out_ctx2;
wire [63:0] MEMC31_burst_count_ctx1;
wire [63:0] MEMC31_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC31(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC31_data_from_Core),
.data_to_Core(MEMC31_data_to_Core),
.valid_ctx1(MEMC31_valid_ctx1),
.addr_out_ctx1(MEMC31_addr_out_ctx1),
.write_en_ctx1(MEMC31_write_en_ctx1),
.start_addr_ctx1(MEMC31_start_addr_ctx1),
.stride_ctx1(MEMC31_stride_ctx1),
.burst_count_ctx1(MEMC31_burst_count_ctx1),
.valid_ctx2(MEMC31_valid_ctx2),
.addr_out_ctx2(MEMC31_addr_out_ctx2),
.write_en_ctx2(MEMC31_write_en_ctx2),
.start_addr_ctx2(MEMC31_start_addr_ctx2),
.stride_ctx2(MEMC31_stride_ctx2),
.burst_count_ctx2(MEMC31_burst_count_ctx2),
.data_in_ctx1(MEMC31_data_in_ctx1),
.data_in_ctx2(MEMC31_data_in_ctx2),
.data_out_ctx1(MEMC31_data_out_ctx1),
.data_out_ctx2(MEMC31_data_out_ctx2),
.write_mem_en_ctx1(MEMC31_write_mem_en_ctx1),
.mem_en_ctx1(MEMC31_mem_en_ctx1),.write_mem_en_ctx2(MEMC31_write_mem_en_ctx2),
.mem_en_ctx2(MEMC31_mem_en_ctx2));

defparam MEMC31.DATA_WIDTH = 32;
defparam MEMC31.ADDR_WIDTH = 6;
defparam MEMC31.STRIDE_WIDTH = 1;
wire MEMC32_valid_ctx1;
wire MEMC32_valid_ctx2;
wire [31:0] MEMC32_data_from_Core;
wire [31:0] MEMC32_data_to_Core;
wire [5:0] MEMC32_addr_out_ctx1;
wire MEMC32_write_en_ctx1;
wire MEMC32_write_mem_en_ctx1;
wire MEMC32_mem_en_ctx1;
wire [5:0] MEMC32_start_addr_ctx1;
wire [0:0] MEMC32_stride_ctx1;
wire [5:0] MEMC32_addr_out_ctx2;
wire MEMC32_write_en_ctx2;
wire MEMC32_write_mem_en_ctx2;
wire MEMC32_mem_en_ctx2;
wire [5:0] MEMC32_start_addr_ctx2;
wire [0:0] MEMC32_stride_ctx2;
wire [31:0] MEMC32_data_in_ctx1;
wire [31:0] MEMC32_data_in_ctx2;
wire [31:0] MEMC32_data_out_ctx1;
wire [31:0] MEMC32_data_out_ctx2;
wire [63:0] MEMC32_burst_count_ctx1;
wire [63:0] MEMC32_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC32(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC32_data_from_Core),
.data_to_Core(MEMC32_data_to_Core),
.valid_ctx1(MEMC32_valid_ctx1),
.addr_out_ctx1(MEMC32_addr_out_ctx1),
.write_en_ctx1(MEMC32_write_en_ctx1),
.start_addr_ctx1(MEMC32_start_addr_ctx1),
.stride_ctx1(MEMC32_stride_ctx1),
.burst_count_ctx1(MEMC32_burst_count_ctx1),
.valid_ctx2(MEMC32_valid_ctx2),
.addr_out_ctx2(MEMC32_addr_out_ctx2),
.write_en_ctx2(MEMC32_write_en_ctx2),
.start_addr_ctx2(MEMC32_start_addr_ctx2),
.stride_ctx2(MEMC32_stride_ctx2),
.burst_count_ctx2(MEMC32_burst_count_ctx2),
.data_in_ctx1(MEMC32_data_in_ctx1),
.data_in_ctx2(MEMC32_data_in_ctx2),
.data_out_ctx1(MEMC32_data_out_ctx1),
.data_out_ctx2(MEMC32_data_out_ctx2),
.write_mem_en_ctx1(MEMC32_write_mem_en_ctx1),
.mem_en_ctx1(MEMC32_mem_en_ctx1),.write_mem_en_ctx2(MEMC32_write_mem_en_ctx2),
.mem_en_ctx2(MEMC32_mem_en_ctx2));

defparam MEMC32.DATA_WIDTH = 32;
defparam MEMC32.ADDR_WIDTH = 6;
defparam MEMC32.STRIDE_WIDTH = 1;
wire MEMC33_valid_ctx1;
wire MEMC33_valid_ctx2;
wire [31:0] MEMC33_data_from_Core;
wire [31:0] MEMC33_data_to_Core;
wire [5:0] MEMC33_addr_out_ctx1;
wire MEMC33_write_en_ctx1;
wire MEMC33_write_mem_en_ctx1;
wire MEMC33_mem_en_ctx1;
wire [5:0] MEMC33_start_addr_ctx1;
wire [0:0] MEMC33_stride_ctx1;
wire [5:0] MEMC33_addr_out_ctx2;
wire MEMC33_write_en_ctx2;
wire MEMC33_write_mem_en_ctx2;
wire MEMC33_mem_en_ctx2;
wire [5:0] MEMC33_start_addr_ctx2;
wire [0:0] MEMC33_stride_ctx2;
wire [31:0] MEMC33_data_in_ctx1;
wire [31:0] MEMC33_data_in_ctx2;
wire [31:0] MEMC33_data_out_ctx1;
wire [31:0] MEMC33_data_out_ctx2;
wire [63:0] MEMC33_burst_count_ctx1;
wire [63:0] MEMC33_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC33(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC33_data_from_Core),
.data_to_Core(MEMC33_data_to_Core),
.valid_ctx1(MEMC33_valid_ctx1),
.addr_out_ctx1(MEMC33_addr_out_ctx1),
.write_en_ctx1(MEMC33_write_en_ctx1),
.start_addr_ctx1(MEMC33_start_addr_ctx1),
.stride_ctx1(MEMC33_stride_ctx1),
.burst_count_ctx1(MEMC33_burst_count_ctx1),
.valid_ctx2(MEMC33_valid_ctx2),
.addr_out_ctx2(MEMC33_addr_out_ctx2),
.write_en_ctx2(MEMC33_write_en_ctx2),
.start_addr_ctx2(MEMC33_start_addr_ctx2),
.stride_ctx2(MEMC33_stride_ctx2),
.burst_count_ctx2(MEMC33_burst_count_ctx2),
.data_in_ctx1(MEMC33_data_in_ctx1),
.data_in_ctx2(MEMC33_data_in_ctx2),
.data_out_ctx1(MEMC33_data_out_ctx1),
.data_out_ctx2(MEMC33_data_out_ctx2),
.write_mem_en_ctx1(MEMC33_write_mem_en_ctx1),
.mem_en_ctx1(MEMC33_mem_en_ctx1),.write_mem_en_ctx2(MEMC33_write_mem_en_ctx2),
.mem_en_ctx2(MEMC33_mem_en_ctx2));

defparam MEMC33.DATA_WIDTH = 32;
defparam MEMC33.ADDR_WIDTH = 6;
defparam MEMC33.STRIDE_WIDTH = 1;
wire MEMC34_valid_ctx1;
wire MEMC34_valid_ctx2;
wire [31:0] MEMC34_data_from_Core;
wire [31:0] MEMC34_data_to_Core;
wire [5:0] MEMC34_addr_out_ctx1;
wire MEMC34_write_en_ctx1;
wire MEMC34_write_mem_en_ctx1;
wire MEMC34_mem_en_ctx1;
wire [5:0] MEMC34_start_addr_ctx1;
wire [0:0] MEMC34_stride_ctx1;
wire [5:0] MEMC34_addr_out_ctx2;
wire MEMC34_write_en_ctx2;
wire MEMC34_write_mem_en_ctx2;
wire MEMC34_mem_en_ctx2;
wire [5:0] MEMC34_start_addr_ctx2;
wire [0:0] MEMC34_stride_ctx2;
wire [31:0] MEMC34_data_in_ctx1;
wire [31:0] MEMC34_data_in_ctx2;
wire [31:0] MEMC34_data_out_ctx1;
wire [31:0] MEMC34_data_out_ctx2;
wire [63:0] MEMC34_burst_count_ctx1;
wire [63:0] MEMC34_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC34(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC34_data_from_Core),
.data_to_Core(MEMC34_data_to_Core),
.valid_ctx1(MEMC34_valid_ctx1),
.addr_out_ctx1(MEMC34_addr_out_ctx1),
.write_en_ctx1(MEMC34_write_en_ctx1),
.start_addr_ctx1(MEMC34_start_addr_ctx1),
.stride_ctx1(MEMC34_stride_ctx1),
.burst_count_ctx1(MEMC34_burst_count_ctx1),
.valid_ctx2(MEMC34_valid_ctx2),
.addr_out_ctx2(MEMC34_addr_out_ctx2),
.write_en_ctx2(MEMC34_write_en_ctx2),
.start_addr_ctx2(MEMC34_start_addr_ctx2),
.stride_ctx2(MEMC34_stride_ctx2),
.burst_count_ctx2(MEMC34_burst_count_ctx2),
.data_in_ctx1(MEMC34_data_in_ctx1),
.data_in_ctx2(MEMC34_data_in_ctx2),
.data_out_ctx1(MEMC34_data_out_ctx1),
.data_out_ctx2(MEMC34_data_out_ctx2),
.write_mem_en_ctx1(MEMC34_write_mem_en_ctx1),
.mem_en_ctx1(MEMC34_mem_en_ctx1),.write_mem_en_ctx2(MEMC34_write_mem_en_ctx2),
.mem_en_ctx2(MEMC34_mem_en_ctx2));

defparam MEMC34.DATA_WIDTH = 32;
defparam MEMC34.ADDR_WIDTH = 6;
defparam MEMC34.STRIDE_WIDTH = 1;
wire MEMC35_valid_ctx1;
wire MEMC35_valid_ctx2;
wire [31:0] MEMC35_data_from_Core;
wire [31:0] MEMC35_data_to_Core;
wire [5:0] MEMC35_addr_out_ctx1;
wire MEMC35_write_en_ctx1;
wire MEMC35_write_mem_en_ctx1;
wire MEMC35_mem_en_ctx1;
wire [5:0] MEMC35_start_addr_ctx1;
wire [0:0] MEMC35_stride_ctx1;
wire [5:0] MEMC35_addr_out_ctx2;
wire MEMC35_write_en_ctx2;
wire MEMC35_write_mem_en_ctx2;
wire MEMC35_mem_en_ctx2;
wire [5:0] MEMC35_start_addr_ctx2;
wire [0:0] MEMC35_stride_ctx2;
wire [31:0] MEMC35_data_in_ctx1;
wire [31:0] MEMC35_data_in_ctx2;
wire [31:0] MEMC35_data_out_ctx1;
wire [31:0] MEMC35_data_out_ctx2;
wire [63:0] MEMC35_burst_count_ctx1;
wire [63:0] MEMC35_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC35(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC35_data_from_Core),
.data_to_Core(MEMC35_data_to_Core),
.valid_ctx1(MEMC35_valid_ctx1),
.addr_out_ctx1(MEMC35_addr_out_ctx1),
.write_en_ctx1(MEMC35_write_en_ctx1),
.start_addr_ctx1(MEMC35_start_addr_ctx1),
.stride_ctx1(MEMC35_stride_ctx1),
.burst_count_ctx1(MEMC35_burst_count_ctx1),
.valid_ctx2(MEMC35_valid_ctx2),
.addr_out_ctx2(MEMC35_addr_out_ctx2),
.write_en_ctx2(MEMC35_write_en_ctx2),
.start_addr_ctx2(MEMC35_start_addr_ctx2),
.stride_ctx2(MEMC35_stride_ctx2),
.burst_count_ctx2(MEMC35_burst_count_ctx2),
.data_in_ctx1(MEMC35_data_in_ctx1),
.data_in_ctx2(MEMC35_data_in_ctx2),
.data_out_ctx1(MEMC35_data_out_ctx1),
.data_out_ctx2(MEMC35_data_out_ctx2),
.write_mem_en_ctx1(MEMC35_write_mem_en_ctx1),
.mem_en_ctx1(MEMC35_mem_en_ctx1),.write_mem_en_ctx2(MEMC35_write_mem_en_ctx2),
.mem_en_ctx2(MEMC35_mem_en_ctx2));

defparam MEMC35.DATA_WIDTH = 32;
defparam MEMC35.ADDR_WIDTH = 6;
defparam MEMC35.STRIDE_WIDTH = 1;
wire MEMC36_valid_ctx1;
wire MEMC36_valid_ctx2;
wire [31:0] MEMC36_data_from_Core;
wire [31:0] MEMC36_data_to_Core;
wire [5:0] MEMC36_addr_out_ctx1;
wire MEMC36_write_en_ctx1;
wire MEMC36_write_mem_en_ctx1;
wire MEMC36_mem_en_ctx1;
wire [5:0] MEMC36_start_addr_ctx1;
wire [0:0] MEMC36_stride_ctx1;
wire [5:0] MEMC36_addr_out_ctx2;
wire MEMC36_write_en_ctx2;
wire MEMC36_write_mem_en_ctx2;
wire MEMC36_mem_en_ctx2;
wire [5:0] MEMC36_start_addr_ctx2;
wire [0:0] MEMC36_stride_ctx2;
wire [31:0] MEMC36_data_in_ctx1;
wire [31:0] MEMC36_data_in_ctx2;
wire [31:0] MEMC36_data_out_ctx1;
wire [31:0] MEMC36_data_out_ctx2;
wire [63:0] MEMC36_burst_count_ctx1;
wire [63:0] MEMC36_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC36(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC36_data_from_Core),
.data_to_Core(MEMC36_data_to_Core),
.valid_ctx1(MEMC36_valid_ctx1),
.addr_out_ctx1(MEMC36_addr_out_ctx1),
.write_en_ctx1(MEMC36_write_en_ctx1),
.start_addr_ctx1(MEMC36_start_addr_ctx1),
.stride_ctx1(MEMC36_stride_ctx1),
.burst_count_ctx1(MEMC36_burst_count_ctx1),
.valid_ctx2(MEMC36_valid_ctx2),
.addr_out_ctx2(MEMC36_addr_out_ctx2),
.write_en_ctx2(MEMC36_write_en_ctx2),
.start_addr_ctx2(MEMC36_start_addr_ctx2),
.stride_ctx2(MEMC36_stride_ctx2),
.burst_count_ctx2(MEMC36_burst_count_ctx2),
.data_in_ctx1(MEMC36_data_in_ctx1),
.data_in_ctx2(MEMC36_data_in_ctx2),
.data_out_ctx1(MEMC36_data_out_ctx1),
.data_out_ctx2(MEMC36_data_out_ctx2),
.write_mem_en_ctx1(MEMC36_write_mem_en_ctx1),
.mem_en_ctx1(MEMC36_mem_en_ctx1),.write_mem_en_ctx2(MEMC36_write_mem_en_ctx2),
.mem_en_ctx2(MEMC36_mem_en_ctx2));

defparam MEMC36.DATA_WIDTH = 32;
defparam MEMC36.ADDR_WIDTH = 6;
defparam MEMC36.STRIDE_WIDTH = 1;
wire MEMC37_valid_ctx1;
wire MEMC37_valid_ctx2;
wire [31:0] MEMC37_data_from_Core;
wire [31:0] MEMC37_data_to_Core;
wire [5:0] MEMC37_addr_out_ctx1;
wire MEMC37_write_en_ctx1;
wire MEMC37_write_mem_en_ctx1;
wire MEMC37_mem_en_ctx1;
wire [5:0] MEMC37_start_addr_ctx1;
wire [0:0] MEMC37_stride_ctx1;
wire [5:0] MEMC37_addr_out_ctx2;
wire MEMC37_write_en_ctx2;
wire MEMC37_write_mem_en_ctx2;
wire MEMC37_mem_en_ctx2;
wire [5:0] MEMC37_start_addr_ctx2;
wire [0:0] MEMC37_stride_ctx2;
wire [31:0] MEMC37_data_in_ctx1;
wire [31:0] MEMC37_data_in_ctx2;
wire [31:0] MEMC37_data_out_ctx1;
wire [31:0] MEMC37_data_out_ctx2;
wire [63:0] MEMC37_burst_count_ctx1;
wire [63:0] MEMC37_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC37(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC37_data_from_Core),
.data_to_Core(MEMC37_data_to_Core),
.valid_ctx1(MEMC37_valid_ctx1),
.addr_out_ctx1(MEMC37_addr_out_ctx1),
.write_en_ctx1(MEMC37_write_en_ctx1),
.start_addr_ctx1(MEMC37_start_addr_ctx1),
.stride_ctx1(MEMC37_stride_ctx1),
.burst_count_ctx1(MEMC37_burst_count_ctx1),
.valid_ctx2(MEMC37_valid_ctx2),
.addr_out_ctx2(MEMC37_addr_out_ctx2),
.write_en_ctx2(MEMC37_write_en_ctx2),
.start_addr_ctx2(MEMC37_start_addr_ctx2),
.stride_ctx2(MEMC37_stride_ctx2),
.burst_count_ctx2(MEMC37_burst_count_ctx2),
.data_in_ctx1(MEMC37_data_in_ctx1),
.data_in_ctx2(MEMC37_data_in_ctx2),
.data_out_ctx1(MEMC37_data_out_ctx1),
.data_out_ctx2(MEMC37_data_out_ctx2),
.write_mem_en_ctx1(MEMC37_write_mem_en_ctx1),
.mem_en_ctx1(MEMC37_mem_en_ctx1),.write_mem_en_ctx2(MEMC37_write_mem_en_ctx2),
.mem_en_ctx2(MEMC37_mem_en_ctx2));

defparam MEMC37.DATA_WIDTH = 32;
defparam MEMC37.ADDR_WIDTH = 6;
defparam MEMC37.STRIDE_WIDTH = 1;
wire MEMC38_valid_ctx1;
wire MEMC38_valid_ctx2;
wire [31:0] MEMC38_data_from_Core;
wire [31:0] MEMC38_data_to_Core;
wire [5:0] MEMC38_addr_out_ctx1;
wire MEMC38_write_en_ctx1;
wire MEMC38_write_mem_en_ctx1;
wire MEMC38_mem_en_ctx1;
wire [5:0] MEMC38_start_addr_ctx1;
wire [0:0] MEMC38_stride_ctx1;
wire [5:0] MEMC38_addr_out_ctx2;
wire MEMC38_write_en_ctx2;
wire MEMC38_write_mem_en_ctx2;
wire MEMC38_mem_en_ctx2;
wire [5:0] MEMC38_start_addr_ctx2;
wire [0:0] MEMC38_stride_ctx2;
wire [31:0] MEMC38_data_in_ctx1;
wire [31:0] MEMC38_data_in_ctx2;
wire [31:0] MEMC38_data_out_ctx1;
wire [31:0] MEMC38_data_out_ctx2;
wire [63:0] MEMC38_burst_count_ctx1;
wire [63:0] MEMC38_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC38(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC38_data_from_Core),
.data_to_Core(MEMC38_data_to_Core),
.valid_ctx1(MEMC38_valid_ctx1),
.addr_out_ctx1(MEMC38_addr_out_ctx1),
.write_en_ctx1(MEMC38_write_en_ctx1),
.start_addr_ctx1(MEMC38_start_addr_ctx1),
.stride_ctx1(MEMC38_stride_ctx1),
.burst_count_ctx1(MEMC38_burst_count_ctx1),
.valid_ctx2(MEMC38_valid_ctx2),
.addr_out_ctx2(MEMC38_addr_out_ctx2),
.write_en_ctx2(MEMC38_write_en_ctx2),
.start_addr_ctx2(MEMC38_start_addr_ctx2),
.stride_ctx2(MEMC38_stride_ctx2),
.burst_count_ctx2(MEMC38_burst_count_ctx2),
.data_in_ctx1(MEMC38_data_in_ctx1),
.data_in_ctx2(MEMC38_data_in_ctx2),
.data_out_ctx1(MEMC38_data_out_ctx1),
.data_out_ctx2(MEMC38_data_out_ctx2),
.write_mem_en_ctx1(MEMC38_write_mem_en_ctx1),
.mem_en_ctx1(MEMC38_mem_en_ctx1),.write_mem_en_ctx2(MEMC38_write_mem_en_ctx2),
.mem_en_ctx2(MEMC38_mem_en_ctx2));

defparam MEMC38.DATA_WIDTH = 32;
defparam MEMC38.ADDR_WIDTH = 6;
defparam MEMC38.STRIDE_WIDTH = 1;
wire MEMC39_valid_ctx1;
wire MEMC39_valid_ctx2;
wire [31:0] MEMC39_data_from_Core;
wire [31:0] MEMC39_data_to_Core;
wire [5:0] MEMC39_addr_out_ctx1;
wire MEMC39_write_en_ctx1;
wire MEMC39_write_mem_en_ctx1;
wire MEMC39_mem_en_ctx1;
wire [5:0] MEMC39_start_addr_ctx1;
wire [0:0] MEMC39_stride_ctx1;
wire [5:0] MEMC39_addr_out_ctx2;
wire MEMC39_write_en_ctx2;
wire MEMC39_write_mem_en_ctx2;
wire MEMC39_mem_en_ctx2;
wire [5:0] MEMC39_start_addr_ctx2;
wire [0:0] MEMC39_stride_ctx2;
wire [31:0] MEMC39_data_in_ctx1;
wire [31:0] MEMC39_data_in_ctx2;
wire [31:0] MEMC39_data_out_ctx1;
wire [31:0] MEMC39_data_out_ctx2;
wire [63:0] MEMC39_burst_count_ctx1;
wire [63:0] MEMC39_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC39(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC39_data_from_Core),
.data_to_Core(MEMC39_data_to_Core),
.valid_ctx1(MEMC39_valid_ctx1),
.addr_out_ctx1(MEMC39_addr_out_ctx1),
.write_en_ctx1(MEMC39_write_en_ctx1),
.start_addr_ctx1(MEMC39_start_addr_ctx1),
.stride_ctx1(MEMC39_stride_ctx1),
.burst_count_ctx1(MEMC39_burst_count_ctx1),
.valid_ctx2(MEMC39_valid_ctx2),
.addr_out_ctx2(MEMC39_addr_out_ctx2),
.write_en_ctx2(MEMC39_write_en_ctx2),
.start_addr_ctx2(MEMC39_start_addr_ctx2),
.stride_ctx2(MEMC39_stride_ctx2),
.burst_count_ctx2(MEMC39_burst_count_ctx2),
.data_in_ctx1(MEMC39_data_in_ctx1),
.data_in_ctx2(MEMC39_data_in_ctx2),
.data_out_ctx1(MEMC39_data_out_ctx1),
.data_out_ctx2(MEMC39_data_out_ctx2),
.write_mem_en_ctx1(MEMC39_write_mem_en_ctx1),
.mem_en_ctx1(MEMC39_mem_en_ctx1),.write_mem_en_ctx2(MEMC39_write_mem_en_ctx2),
.mem_en_ctx2(MEMC39_mem_en_ctx2));

defparam MEMC39.DATA_WIDTH = 32;
defparam MEMC39.ADDR_WIDTH = 6;
defparam MEMC39.STRIDE_WIDTH = 1;
wire MEMC40_valid_ctx1;
wire MEMC40_valid_ctx2;
wire [31:0] MEMC40_data_from_Core;
wire [31:0] MEMC40_data_to_Core;
wire [5:0] MEMC40_addr_out_ctx1;
wire MEMC40_write_en_ctx1;
wire MEMC40_write_mem_en_ctx1;
wire MEMC40_mem_en_ctx1;
wire [5:0] MEMC40_start_addr_ctx1;
wire [0:0] MEMC40_stride_ctx1;
wire [5:0] MEMC40_addr_out_ctx2;
wire MEMC40_write_en_ctx2;
wire MEMC40_write_mem_en_ctx2;
wire MEMC40_mem_en_ctx2;
wire [5:0] MEMC40_start_addr_ctx2;
wire [0:0] MEMC40_stride_ctx2;
wire [31:0] MEMC40_data_in_ctx1;
wire [31:0] MEMC40_data_in_ctx2;
wire [31:0] MEMC40_data_out_ctx1;
wire [31:0] MEMC40_data_out_ctx2;
wire [63:0] MEMC40_burst_count_ctx1;
wire [63:0] MEMC40_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC40(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC40_data_from_Core),
.data_to_Core(MEMC40_data_to_Core),
.valid_ctx1(MEMC40_valid_ctx1),
.addr_out_ctx1(MEMC40_addr_out_ctx1),
.write_en_ctx1(MEMC40_write_en_ctx1),
.start_addr_ctx1(MEMC40_start_addr_ctx1),
.stride_ctx1(MEMC40_stride_ctx1),
.burst_count_ctx1(MEMC40_burst_count_ctx1),
.valid_ctx2(MEMC40_valid_ctx2),
.addr_out_ctx2(MEMC40_addr_out_ctx2),
.write_en_ctx2(MEMC40_write_en_ctx2),
.start_addr_ctx2(MEMC40_start_addr_ctx2),
.stride_ctx2(MEMC40_stride_ctx2),
.burst_count_ctx2(MEMC40_burst_count_ctx2),
.data_in_ctx1(MEMC40_data_in_ctx1),
.data_in_ctx2(MEMC40_data_in_ctx2),
.data_out_ctx1(MEMC40_data_out_ctx1),
.data_out_ctx2(MEMC40_data_out_ctx2),
.write_mem_en_ctx1(MEMC40_write_mem_en_ctx1),
.mem_en_ctx1(MEMC40_mem_en_ctx1),.write_mem_en_ctx2(MEMC40_write_mem_en_ctx2),
.mem_en_ctx2(MEMC40_mem_en_ctx2));

defparam MEMC40.DATA_WIDTH = 32;
defparam MEMC40.ADDR_WIDTH = 6;
defparam MEMC40.STRIDE_WIDTH = 1;
wire MEMC41_valid_ctx1;
wire MEMC41_valid_ctx2;
wire [31:0] MEMC41_data_from_Core;
wire [31:0] MEMC41_data_to_Core;
wire [5:0] MEMC41_addr_out_ctx1;
wire MEMC41_write_en_ctx1;
wire MEMC41_write_mem_en_ctx1;
wire MEMC41_mem_en_ctx1;
wire [5:0] MEMC41_start_addr_ctx1;
wire [0:0] MEMC41_stride_ctx1;
wire [5:0] MEMC41_addr_out_ctx2;
wire MEMC41_write_en_ctx2;
wire MEMC41_write_mem_en_ctx2;
wire MEMC41_mem_en_ctx2;
wire [5:0] MEMC41_start_addr_ctx2;
wire [0:0] MEMC41_stride_ctx2;
wire [31:0] MEMC41_data_in_ctx1;
wire [31:0] MEMC41_data_in_ctx2;
wire [31:0] MEMC41_data_out_ctx1;
wire [31:0] MEMC41_data_out_ctx2;
wire [63:0] MEMC41_burst_count_ctx1;
wire [63:0] MEMC41_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC41(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC41_data_from_Core),
.data_to_Core(MEMC41_data_to_Core),
.valid_ctx1(MEMC41_valid_ctx1),
.addr_out_ctx1(MEMC41_addr_out_ctx1),
.write_en_ctx1(MEMC41_write_en_ctx1),
.start_addr_ctx1(MEMC41_start_addr_ctx1),
.stride_ctx1(MEMC41_stride_ctx1),
.burst_count_ctx1(MEMC41_burst_count_ctx1),
.valid_ctx2(MEMC41_valid_ctx2),
.addr_out_ctx2(MEMC41_addr_out_ctx2),
.write_en_ctx2(MEMC41_write_en_ctx2),
.start_addr_ctx2(MEMC41_start_addr_ctx2),
.stride_ctx2(MEMC41_stride_ctx2),
.burst_count_ctx2(MEMC41_burst_count_ctx2),
.data_in_ctx1(MEMC41_data_in_ctx1),
.data_in_ctx2(MEMC41_data_in_ctx2),
.data_out_ctx1(MEMC41_data_out_ctx1),
.data_out_ctx2(MEMC41_data_out_ctx2),
.write_mem_en_ctx1(MEMC41_write_mem_en_ctx1),
.mem_en_ctx1(MEMC41_mem_en_ctx1),.write_mem_en_ctx2(MEMC41_write_mem_en_ctx2),
.mem_en_ctx2(MEMC41_mem_en_ctx2));

defparam MEMC41.DATA_WIDTH = 32;
defparam MEMC41.ADDR_WIDTH = 6;
defparam MEMC41.STRIDE_WIDTH = 1;
wire MEMC42_valid_ctx1;
wire MEMC42_valid_ctx2;
wire [31:0] MEMC42_data_from_Core;
wire [31:0] MEMC42_data_to_Core;
wire [5:0] MEMC42_addr_out_ctx1;
wire MEMC42_write_en_ctx1;
wire MEMC42_write_mem_en_ctx1;
wire MEMC42_mem_en_ctx1;
wire [5:0] MEMC42_start_addr_ctx1;
wire [0:0] MEMC42_stride_ctx1;
wire [5:0] MEMC42_addr_out_ctx2;
wire MEMC42_write_en_ctx2;
wire MEMC42_write_mem_en_ctx2;
wire MEMC42_mem_en_ctx2;
wire [5:0] MEMC42_start_addr_ctx2;
wire [0:0] MEMC42_stride_ctx2;
wire [31:0] MEMC42_data_in_ctx1;
wire [31:0] MEMC42_data_in_ctx2;
wire [31:0] MEMC42_data_out_ctx1;
wire [31:0] MEMC42_data_out_ctx2;
wire [63:0] MEMC42_burst_count_ctx1;
wire [63:0] MEMC42_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC42(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC42_data_from_Core),
.data_to_Core(MEMC42_data_to_Core),
.valid_ctx1(MEMC42_valid_ctx1),
.addr_out_ctx1(MEMC42_addr_out_ctx1),
.write_en_ctx1(MEMC42_write_en_ctx1),
.start_addr_ctx1(MEMC42_start_addr_ctx1),
.stride_ctx1(MEMC42_stride_ctx1),
.burst_count_ctx1(MEMC42_burst_count_ctx1),
.valid_ctx2(MEMC42_valid_ctx2),
.addr_out_ctx2(MEMC42_addr_out_ctx2),
.write_en_ctx2(MEMC42_write_en_ctx2),
.start_addr_ctx2(MEMC42_start_addr_ctx2),
.stride_ctx2(MEMC42_stride_ctx2),
.burst_count_ctx2(MEMC42_burst_count_ctx2),
.data_in_ctx1(MEMC42_data_in_ctx1),
.data_in_ctx2(MEMC42_data_in_ctx2),
.data_out_ctx1(MEMC42_data_out_ctx1),
.data_out_ctx2(MEMC42_data_out_ctx2),
.write_mem_en_ctx1(MEMC42_write_mem_en_ctx1),
.mem_en_ctx1(MEMC42_mem_en_ctx1),.write_mem_en_ctx2(MEMC42_write_mem_en_ctx2),
.mem_en_ctx2(MEMC42_mem_en_ctx2));

defparam MEMC42.DATA_WIDTH = 32;
defparam MEMC42.ADDR_WIDTH = 6;
defparam MEMC42.STRIDE_WIDTH = 1;
wire MEMC43_valid_ctx1;
wire MEMC43_valid_ctx2;
wire [31:0] MEMC43_data_from_Core;
wire [31:0] MEMC43_data_to_Core;
wire [5:0] MEMC43_addr_out_ctx1;
wire MEMC43_write_en_ctx1;
wire MEMC43_write_mem_en_ctx1;
wire MEMC43_mem_en_ctx1;
wire [5:0] MEMC43_start_addr_ctx1;
wire [0:0] MEMC43_stride_ctx1;
wire [5:0] MEMC43_addr_out_ctx2;
wire MEMC43_write_en_ctx2;
wire MEMC43_write_mem_en_ctx2;
wire MEMC43_mem_en_ctx2;
wire [5:0] MEMC43_start_addr_ctx2;
wire [0:0] MEMC43_stride_ctx2;
wire [31:0] MEMC43_data_in_ctx1;
wire [31:0] MEMC43_data_in_ctx2;
wire [31:0] MEMC43_data_out_ctx1;
wire [31:0] MEMC43_data_out_ctx2;
wire [63:0] MEMC43_burst_count_ctx1;
wire [63:0] MEMC43_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC43(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC43_data_from_Core),
.data_to_Core(MEMC43_data_to_Core),
.valid_ctx1(MEMC43_valid_ctx1),
.addr_out_ctx1(MEMC43_addr_out_ctx1),
.write_en_ctx1(MEMC43_write_en_ctx1),
.start_addr_ctx1(MEMC43_start_addr_ctx1),
.stride_ctx1(MEMC43_stride_ctx1),
.burst_count_ctx1(MEMC43_burst_count_ctx1),
.valid_ctx2(MEMC43_valid_ctx2),
.addr_out_ctx2(MEMC43_addr_out_ctx2),
.write_en_ctx2(MEMC43_write_en_ctx2),
.start_addr_ctx2(MEMC43_start_addr_ctx2),
.stride_ctx2(MEMC43_stride_ctx2),
.burst_count_ctx2(MEMC43_burst_count_ctx2),
.data_in_ctx1(MEMC43_data_in_ctx1),
.data_in_ctx2(MEMC43_data_in_ctx2),
.data_out_ctx1(MEMC43_data_out_ctx1),
.data_out_ctx2(MEMC43_data_out_ctx2),
.write_mem_en_ctx1(MEMC43_write_mem_en_ctx1),
.mem_en_ctx1(MEMC43_mem_en_ctx1),.write_mem_en_ctx2(MEMC43_write_mem_en_ctx2),
.mem_en_ctx2(MEMC43_mem_en_ctx2));

defparam MEMC43.DATA_WIDTH = 32;
defparam MEMC43.ADDR_WIDTH = 6;
defparam MEMC43.STRIDE_WIDTH = 1;
wire MEMC44_valid_ctx1;
wire MEMC44_valid_ctx2;
wire [31:0] MEMC44_data_from_Core;
wire [31:0] MEMC44_data_to_Core;
wire [5:0] MEMC44_addr_out_ctx1;
wire MEMC44_write_en_ctx1;
wire MEMC44_write_mem_en_ctx1;
wire MEMC44_mem_en_ctx1;
wire [5:0] MEMC44_start_addr_ctx1;
wire [0:0] MEMC44_stride_ctx1;
wire [5:0] MEMC44_addr_out_ctx2;
wire MEMC44_write_en_ctx2;
wire MEMC44_write_mem_en_ctx2;
wire MEMC44_mem_en_ctx2;
wire [5:0] MEMC44_start_addr_ctx2;
wire [0:0] MEMC44_stride_ctx2;
wire [31:0] MEMC44_data_in_ctx1;
wire [31:0] MEMC44_data_in_ctx2;
wire [31:0] MEMC44_data_out_ctx1;
wire [31:0] MEMC44_data_out_ctx2;
wire [63:0] MEMC44_burst_count_ctx1;
wire [63:0] MEMC44_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC44(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC44_data_from_Core),
.data_to_Core(MEMC44_data_to_Core),
.valid_ctx1(MEMC44_valid_ctx1),
.addr_out_ctx1(MEMC44_addr_out_ctx1),
.write_en_ctx1(MEMC44_write_en_ctx1),
.start_addr_ctx1(MEMC44_start_addr_ctx1),
.stride_ctx1(MEMC44_stride_ctx1),
.burst_count_ctx1(MEMC44_burst_count_ctx1),
.valid_ctx2(MEMC44_valid_ctx2),
.addr_out_ctx2(MEMC44_addr_out_ctx2),
.write_en_ctx2(MEMC44_write_en_ctx2),
.start_addr_ctx2(MEMC44_start_addr_ctx2),
.stride_ctx2(MEMC44_stride_ctx2),
.burst_count_ctx2(MEMC44_burst_count_ctx2),
.data_in_ctx1(MEMC44_data_in_ctx1),
.data_in_ctx2(MEMC44_data_in_ctx2),
.data_out_ctx1(MEMC44_data_out_ctx1),
.data_out_ctx2(MEMC44_data_out_ctx2),
.write_mem_en_ctx1(MEMC44_write_mem_en_ctx1),
.mem_en_ctx1(MEMC44_mem_en_ctx1),.write_mem_en_ctx2(MEMC44_write_mem_en_ctx2),
.mem_en_ctx2(MEMC44_mem_en_ctx2));

defparam MEMC44.DATA_WIDTH = 32;
defparam MEMC44.ADDR_WIDTH = 6;
defparam MEMC44.STRIDE_WIDTH = 1;
wire MEMC45_valid_ctx1;
wire MEMC45_valid_ctx2;
wire [31:0] MEMC45_data_from_Core;
wire [31:0] MEMC45_data_to_Core;
wire [5:0] MEMC45_addr_out_ctx1;
wire MEMC45_write_en_ctx1;
wire MEMC45_write_mem_en_ctx1;
wire MEMC45_mem_en_ctx1;
wire [5:0] MEMC45_start_addr_ctx1;
wire [0:0] MEMC45_stride_ctx1;
wire [5:0] MEMC45_addr_out_ctx2;
wire MEMC45_write_en_ctx2;
wire MEMC45_write_mem_en_ctx2;
wire MEMC45_mem_en_ctx2;
wire [5:0] MEMC45_start_addr_ctx2;
wire [0:0] MEMC45_stride_ctx2;
wire [31:0] MEMC45_data_in_ctx1;
wire [31:0] MEMC45_data_in_ctx2;
wire [31:0] MEMC45_data_out_ctx1;
wire [31:0] MEMC45_data_out_ctx2;
wire [63:0] MEMC45_burst_count_ctx1;
wire [63:0] MEMC45_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC45(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC45_data_from_Core),
.data_to_Core(MEMC45_data_to_Core),
.valid_ctx1(MEMC45_valid_ctx1),
.addr_out_ctx1(MEMC45_addr_out_ctx1),
.write_en_ctx1(MEMC45_write_en_ctx1),
.start_addr_ctx1(MEMC45_start_addr_ctx1),
.stride_ctx1(MEMC45_stride_ctx1),
.burst_count_ctx1(MEMC45_burst_count_ctx1),
.valid_ctx2(MEMC45_valid_ctx2),
.addr_out_ctx2(MEMC45_addr_out_ctx2),
.write_en_ctx2(MEMC45_write_en_ctx2),
.start_addr_ctx2(MEMC45_start_addr_ctx2),
.stride_ctx2(MEMC45_stride_ctx2),
.burst_count_ctx2(MEMC45_burst_count_ctx2),
.data_in_ctx1(MEMC45_data_in_ctx1),
.data_in_ctx2(MEMC45_data_in_ctx2),
.data_out_ctx1(MEMC45_data_out_ctx1),
.data_out_ctx2(MEMC45_data_out_ctx2),
.write_mem_en_ctx1(MEMC45_write_mem_en_ctx1),
.mem_en_ctx1(MEMC45_mem_en_ctx1),.write_mem_en_ctx2(MEMC45_write_mem_en_ctx2),
.mem_en_ctx2(MEMC45_mem_en_ctx2));

defparam MEMC45.DATA_WIDTH = 32;
defparam MEMC45.ADDR_WIDTH = 6;
defparam MEMC45.STRIDE_WIDTH = 1;
wire MEMC46_valid_ctx1;
wire MEMC46_valid_ctx2;
wire [31:0] MEMC46_data_from_Core;
wire [31:0] MEMC46_data_to_Core;
wire [5:0] MEMC46_addr_out_ctx1;
wire MEMC46_write_en_ctx1;
wire MEMC46_write_mem_en_ctx1;
wire MEMC46_mem_en_ctx1;
wire [5:0] MEMC46_start_addr_ctx1;
wire [0:0] MEMC46_stride_ctx1;
wire [5:0] MEMC46_addr_out_ctx2;
wire MEMC46_write_en_ctx2;
wire MEMC46_write_mem_en_ctx2;
wire MEMC46_mem_en_ctx2;
wire [5:0] MEMC46_start_addr_ctx2;
wire [0:0] MEMC46_stride_ctx2;
wire [31:0] MEMC46_data_in_ctx1;
wire [31:0] MEMC46_data_in_ctx2;
wire [31:0] MEMC46_data_out_ctx1;
wire [31:0] MEMC46_data_out_ctx2;
wire [63:0] MEMC46_burst_count_ctx1;
wire [63:0] MEMC46_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC46(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC46_data_from_Core),
.data_to_Core(MEMC46_data_to_Core),
.valid_ctx1(MEMC46_valid_ctx1),
.addr_out_ctx1(MEMC46_addr_out_ctx1),
.write_en_ctx1(MEMC46_write_en_ctx1),
.start_addr_ctx1(MEMC46_start_addr_ctx1),
.stride_ctx1(MEMC46_stride_ctx1),
.burst_count_ctx1(MEMC46_burst_count_ctx1),
.valid_ctx2(MEMC46_valid_ctx2),
.addr_out_ctx2(MEMC46_addr_out_ctx2),
.write_en_ctx2(MEMC46_write_en_ctx2),
.start_addr_ctx2(MEMC46_start_addr_ctx2),
.stride_ctx2(MEMC46_stride_ctx2),
.burst_count_ctx2(MEMC46_burst_count_ctx2),
.data_in_ctx1(MEMC46_data_in_ctx1),
.data_in_ctx2(MEMC46_data_in_ctx2),
.data_out_ctx1(MEMC46_data_out_ctx1),
.data_out_ctx2(MEMC46_data_out_ctx2),
.write_mem_en_ctx1(MEMC46_write_mem_en_ctx1),
.mem_en_ctx1(MEMC46_mem_en_ctx1),.write_mem_en_ctx2(MEMC46_write_mem_en_ctx2),
.mem_en_ctx2(MEMC46_mem_en_ctx2));

defparam MEMC46.DATA_WIDTH = 32;
defparam MEMC46.ADDR_WIDTH = 6;
defparam MEMC46.STRIDE_WIDTH = 1;
wire MEMC47_valid_ctx1;
wire MEMC47_valid_ctx2;
wire [31:0] MEMC47_data_from_Core;
wire [31:0] MEMC47_data_to_Core;
wire [5:0] MEMC47_addr_out_ctx1;
wire MEMC47_write_en_ctx1;
wire MEMC47_write_mem_en_ctx1;
wire MEMC47_mem_en_ctx1;
wire [5:0] MEMC47_start_addr_ctx1;
wire [0:0] MEMC47_stride_ctx1;
wire [5:0] MEMC47_addr_out_ctx2;
wire MEMC47_write_en_ctx2;
wire MEMC47_write_mem_en_ctx2;
wire MEMC47_mem_en_ctx2;
wire [5:0] MEMC47_start_addr_ctx2;
wire [0:0] MEMC47_stride_ctx2;
wire [31:0] MEMC47_data_in_ctx1;
wire [31:0] MEMC47_data_in_ctx2;
wire [31:0] MEMC47_data_out_ctx1;
wire [31:0] MEMC47_data_out_ctx2;
wire [63:0] MEMC47_burst_count_ctx1;
wire [63:0] MEMC47_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC47(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC47_data_from_Core),
.data_to_Core(MEMC47_data_to_Core),
.valid_ctx1(MEMC47_valid_ctx1),
.addr_out_ctx1(MEMC47_addr_out_ctx1),
.write_en_ctx1(MEMC47_write_en_ctx1),
.start_addr_ctx1(MEMC47_start_addr_ctx1),
.stride_ctx1(MEMC47_stride_ctx1),
.burst_count_ctx1(MEMC47_burst_count_ctx1),
.valid_ctx2(MEMC47_valid_ctx2),
.addr_out_ctx2(MEMC47_addr_out_ctx2),
.write_en_ctx2(MEMC47_write_en_ctx2),
.start_addr_ctx2(MEMC47_start_addr_ctx2),
.stride_ctx2(MEMC47_stride_ctx2),
.burst_count_ctx2(MEMC47_burst_count_ctx2),
.data_in_ctx1(MEMC47_data_in_ctx1),
.data_in_ctx2(MEMC47_data_in_ctx2),
.data_out_ctx1(MEMC47_data_out_ctx1),
.data_out_ctx2(MEMC47_data_out_ctx2),
.write_mem_en_ctx1(MEMC47_write_mem_en_ctx1),
.mem_en_ctx1(MEMC47_mem_en_ctx1),.write_mem_en_ctx2(MEMC47_write_mem_en_ctx2),
.mem_en_ctx2(MEMC47_mem_en_ctx2));

defparam MEMC47.DATA_WIDTH = 32;
defparam MEMC47.ADDR_WIDTH = 6;
defparam MEMC47.STRIDE_WIDTH = 1;
wire MEMC48_valid_ctx1;
wire MEMC48_valid_ctx2;
wire [31:0] MEMC48_data_from_Core;
wire [31:0] MEMC48_data_to_Core;
wire [5:0] MEMC48_addr_out_ctx1;
wire MEMC48_write_en_ctx1;
wire MEMC48_write_mem_en_ctx1;
wire MEMC48_mem_en_ctx1;
wire [5:0] MEMC48_start_addr_ctx1;
wire [0:0] MEMC48_stride_ctx1;
wire [5:0] MEMC48_addr_out_ctx2;
wire MEMC48_write_en_ctx2;
wire MEMC48_write_mem_en_ctx2;
wire MEMC48_mem_en_ctx2;
wire [5:0] MEMC48_start_addr_ctx2;
wire [0:0] MEMC48_stride_ctx2;
wire [31:0] MEMC48_data_in_ctx1;
wire [31:0] MEMC48_data_in_ctx2;
wire [31:0] MEMC48_data_out_ctx1;
wire [31:0] MEMC48_data_out_ctx2;
wire [63:0] MEMC48_burst_count_ctx1;
wire [63:0] MEMC48_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC48(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC48_data_from_Core),
.data_to_Core(MEMC48_data_to_Core),
.valid_ctx1(MEMC48_valid_ctx1),
.addr_out_ctx1(MEMC48_addr_out_ctx1),
.write_en_ctx1(MEMC48_write_en_ctx1),
.start_addr_ctx1(MEMC48_start_addr_ctx1),
.stride_ctx1(MEMC48_stride_ctx1),
.burst_count_ctx1(MEMC48_burst_count_ctx1),
.valid_ctx2(MEMC48_valid_ctx2),
.addr_out_ctx2(MEMC48_addr_out_ctx2),
.write_en_ctx2(MEMC48_write_en_ctx2),
.start_addr_ctx2(MEMC48_start_addr_ctx2),
.stride_ctx2(MEMC48_stride_ctx2),
.burst_count_ctx2(MEMC48_burst_count_ctx2),
.data_in_ctx1(MEMC48_data_in_ctx1),
.data_in_ctx2(MEMC48_data_in_ctx2),
.data_out_ctx1(MEMC48_data_out_ctx1),
.data_out_ctx2(MEMC48_data_out_ctx2),
.write_mem_en_ctx1(MEMC48_write_mem_en_ctx1),
.mem_en_ctx1(MEMC48_mem_en_ctx1),.write_mem_en_ctx2(MEMC48_write_mem_en_ctx2),
.mem_en_ctx2(MEMC48_mem_en_ctx2));

defparam MEMC48.DATA_WIDTH = 32;
defparam MEMC48.ADDR_WIDTH = 6;
defparam MEMC48.STRIDE_WIDTH = 1;
wire MEMC49_valid_ctx1;
wire MEMC49_valid_ctx2;
wire [31:0] MEMC49_data_from_Core;
wire [31:0] MEMC49_data_to_Core;
wire [5:0] MEMC49_addr_out_ctx1;
wire MEMC49_write_en_ctx1;
wire MEMC49_write_mem_en_ctx1;
wire MEMC49_mem_en_ctx1;
wire [5:0] MEMC49_start_addr_ctx1;
wire [0:0] MEMC49_stride_ctx1;
wire [5:0] MEMC49_addr_out_ctx2;
wire MEMC49_write_en_ctx2;
wire MEMC49_write_mem_en_ctx2;
wire MEMC49_mem_en_ctx2;
wire [5:0] MEMC49_start_addr_ctx2;
wire [0:0] MEMC49_stride_ctx2;
wire [31:0] MEMC49_data_in_ctx1;
wire [31:0] MEMC49_data_in_ctx2;
wire [31:0] MEMC49_data_out_ctx1;
wire [31:0] MEMC49_data_out_ctx2;
wire [63:0] MEMC49_burst_count_ctx1;
wire [63:0] MEMC49_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC49(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC49_data_from_Core),
.data_to_Core(MEMC49_data_to_Core),
.valid_ctx1(MEMC49_valid_ctx1),
.addr_out_ctx1(MEMC49_addr_out_ctx1),
.write_en_ctx1(MEMC49_write_en_ctx1),
.start_addr_ctx1(MEMC49_start_addr_ctx1),
.stride_ctx1(MEMC49_stride_ctx1),
.burst_count_ctx1(MEMC49_burst_count_ctx1),
.valid_ctx2(MEMC49_valid_ctx2),
.addr_out_ctx2(MEMC49_addr_out_ctx2),
.write_en_ctx2(MEMC49_write_en_ctx2),
.start_addr_ctx2(MEMC49_start_addr_ctx2),
.stride_ctx2(MEMC49_stride_ctx2),
.burst_count_ctx2(MEMC49_burst_count_ctx2),
.data_in_ctx1(MEMC49_data_in_ctx1),
.data_in_ctx2(MEMC49_data_in_ctx2),
.data_out_ctx1(MEMC49_data_out_ctx1),
.data_out_ctx2(MEMC49_data_out_ctx2),
.write_mem_en_ctx1(MEMC49_write_mem_en_ctx1),
.mem_en_ctx1(MEMC49_mem_en_ctx1),.write_mem_en_ctx2(MEMC49_write_mem_en_ctx2),
.mem_en_ctx2(MEMC49_mem_en_ctx2));

defparam MEMC49.DATA_WIDTH = 32;
defparam MEMC49.ADDR_WIDTH = 6;
defparam MEMC49.STRIDE_WIDTH = 1;
wire MEMC50_valid_ctx1;
wire MEMC50_valid_ctx2;
wire [31:0] MEMC50_data_from_Core;
wire [31:0] MEMC50_data_to_Core;
wire [5:0] MEMC50_addr_out_ctx1;
wire MEMC50_write_en_ctx1;
wire MEMC50_write_mem_en_ctx1;
wire MEMC50_mem_en_ctx1;
wire [5:0] MEMC50_start_addr_ctx1;
wire [0:0] MEMC50_stride_ctx1;
wire [5:0] MEMC50_addr_out_ctx2;
wire MEMC50_write_en_ctx2;
wire MEMC50_write_mem_en_ctx2;
wire MEMC50_mem_en_ctx2;
wire [5:0] MEMC50_start_addr_ctx2;
wire [0:0] MEMC50_stride_ctx2;
wire [31:0] MEMC50_data_in_ctx1;
wire [31:0] MEMC50_data_in_ctx2;
wire [31:0] MEMC50_data_out_ctx1;
wire [31:0] MEMC50_data_out_ctx2;
wire [63:0] MEMC50_burst_count_ctx1;
wire [63:0] MEMC50_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC50(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC50_data_from_Core),
.data_to_Core(MEMC50_data_to_Core),
.valid_ctx1(MEMC50_valid_ctx1),
.addr_out_ctx1(MEMC50_addr_out_ctx1),
.write_en_ctx1(MEMC50_write_en_ctx1),
.start_addr_ctx1(MEMC50_start_addr_ctx1),
.stride_ctx1(MEMC50_stride_ctx1),
.burst_count_ctx1(MEMC50_burst_count_ctx1),
.valid_ctx2(MEMC50_valid_ctx2),
.addr_out_ctx2(MEMC50_addr_out_ctx2),
.write_en_ctx2(MEMC50_write_en_ctx2),
.start_addr_ctx2(MEMC50_start_addr_ctx2),
.stride_ctx2(MEMC50_stride_ctx2),
.burst_count_ctx2(MEMC50_burst_count_ctx2),
.data_in_ctx1(MEMC50_data_in_ctx1),
.data_in_ctx2(MEMC50_data_in_ctx2),
.data_out_ctx1(MEMC50_data_out_ctx1),
.data_out_ctx2(MEMC50_data_out_ctx2),
.write_mem_en_ctx1(MEMC50_write_mem_en_ctx1),
.mem_en_ctx1(MEMC50_mem_en_ctx1),.write_mem_en_ctx2(MEMC50_write_mem_en_ctx2),
.mem_en_ctx2(MEMC50_mem_en_ctx2));

defparam MEMC50.DATA_WIDTH = 32;
defparam MEMC50.ADDR_WIDTH = 6;
defparam MEMC50.STRIDE_WIDTH = 1;
wire MEMC51_valid_ctx1;
wire MEMC51_valid_ctx2;
wire [31:0] MEMC51_data_from_Core;
wire [31:0] MEMC51_data_to_Core;
wire [5:0] MEMC51_addr_out_ctx1;
wire MEMC51_write_en_ctx1;
wire MEMC51_write_mem_en_ctx1;
wire MEMC51_mem_en_ctx1;
wire [5:0] MEMC51_start_addr_ctx1;
wire [0:0] MEMC51_stride_ctx1;
wire [5:0] MEMC51_addr_out_ctx2;
wire MEMC51_write_en_ctx2;
wire MEMC51_write_mem_en_ctx2;
wire MEMC51_mem_en_ctx2;
wire [5:0] MEMC51_start_addr_ctx2;
wire [0:0] MEMC51_stride_ctx2;
wire [31:0] MEMC51_data_in_ctx1;
wire [31:0] MEMC51_data_in_ctx2;
wire [31:0] MEMC51_data_out_ctx1;
wire [31:0] MEMC51_data_out_ctx2;
wire [63:0] MEMC51_burst_count_ctx1;
wire [63:0] MEMC51_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC51(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC51_data_from_Core),
.data_to_Core(MEMC51_data_to_Core),
.valid_ctx1(MEMC51_valid_ctx1),
.addr_out_ctx1(MEMC51_addr_out_ctx1),
.write_en_ctx1(MEMC51_write_en_ctx1),
.start_addr_ctx1(MEMC51_start_addr_ctx1),
.stride_ctx1(MEMC51_stride_ctx1),
.burst_count_ctx1(MEMC51_burst_count_ctx1),
.valid_ctx2(MEMC51_valid_ctx2),
.addr_out_ctx2(MEMC51_addr_out_ctx2),
.write_en_ctx2(MEMC51_write_en_ctx2),
.start_addr_ctx2(MEMC51_start_addr_ctx2),
.stride_ctx2(MEMC51_stride_ctx2),
.burst_count_ctx2(MEMC51_burst_count_ctx2),
.data_in_ctx1(MEMC51_data_in_ctx1),
.data_in_ctx2(MEMC51_data_in_ctx2),
.data_out_ctx1(MEMC51_data_out_ctx1),
.data_out_ctx2(MEMC51_data_out_ctx2),
.write_mem_en_ctx1(MEMC51_write_mem_en_ctx1),
.mem_en_ctx1(MEMC51_mem_en_ctx1),.write_mem_en_ctx2(MEMC51_write_mem_en_ctx2),
.mem_en_ctx2(MEMC51_mem_en_ctx2));

defparam MEMC51.DATA_WIDTH = 32;
defparam MEMC51.ADDR_WIDTH = 6;
defparam MEMC51.STRIDE_WIDTH = 1;
wire MEMC52_valid_ctx1;
wire MEMC52_valid_ctx2;
wire [31:0] MEMC52_data_from_Core;
wire [31:0] MEMC52_data_to_Core;
wire [5:0] MEMC52_addr_out_ctx1;
wire MEMC52_write_en_ctx1;
wire MEMC52_write_mem_en_ctx1;
wire MEMC52_mem_en_ctx1;
wire [5:0] MEMC52_start_addr_ctx1;
wire [0:0] MEMC52_stride_ctx1;
wire [5:0] MEMC52_addr_out_ctx2;
wire MEMC52_write_en_ctx2;
wire MEMC52_write_mem_en_ctx2;
wire MEMC52_mem_en_ctx2;
wire [5:0] MEMC52_start_addr_ctx2;
wire [0:0] MEMC52_stride_ctx2;
wire [31:0] MEMC52_data_in_ctx1;
wire [31:0] MEMC52_data_in_ctx2;
wire [31:0] MEMC52_data_out_ctx1;
wire [31:0] MEMC52_data_out_ctx2;
wire [63:0] MEMC52_burst_count_ctx1;
wire [63:0] MEMC52_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC52(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC52_data_from_Core),
.data_to_Core(MEMC52_data_to_Core),
.valid_ctx1(MEMC52_valid_ctx1),
.addr_out_ctx1(MEMC52_addr_out_ctx1),
.write_en_ctx1(MEMC52_write_en_ctx1),
.start_addr_ctx1(MEMC52_start_addr_ctx1),
.stride_ctx1(MEMC52_stride_ctx1),
.burst_count_ctx1(MEMC52_burst_count_ctx1),
.valid_ctx2(MEMC52_valid_ctx2),
.addr_out_ctx2(MEMC52_addr_out_ctx2),
.write_en_ctx2(MEMC52_write_en_ctx2),
.start_addr_ctx2(MEMC52_start_addr_ctx2),
.stride_ctx2(MEMC52_stride_ctx2),
.burst_count_ctx2(MEMC52_burst_count_ctx2),
.data_in_ctx1(MEMC52_data_in_ctx1),
.data_in_ctx2(MEMC52_data_in_ctx2),
.data_out_ctx1(MEMC52_data_out_ctx1),
.data_out_ctx2(MEMC52_data_out_ctx2),
.write_mem_en_ctx1(MEMC52_write_mem_en_ctx1),
.mem_en_ctx1(MEMC52_mem_en_ctx1),.write_mem_en_ctx2(MEMC52_write_mem_en_ctx2),
.mem_en_ctx2(MEMC52_mem_en_ctx2));

defparam MEMC52.DATA_WIDTH = 32;
defparam MEMC52.ADDR_WIDTH = 6;
defparam MEMC52.STRIDE_WIDTH = 1;
wire MEMC53_valid_ctx1;
wire MEMC53_valid_ctx2;
wire [31:0] MEMC53_data_from_Core;
wire [31:0] MEMC53_data_to_Core;
wire [5:0] MEMC53_addr_out_ctx1;
wire MEMC53_write_en_ctx1;
wire MEMC53_write_mem_en_ctx1;
wire MEMC53_mem_en_ctx1;
wire [5:0] MEMC53_start_addr_ctx1;
wire [0:0] MEMC53_stride_ctx1;
wire [5:0] MEMC53_addr_out_ctx2;
wire MEMC53_write_en_ctx2;
wire MEMC53_write_mem_en_ctx2;
wire MEMC53_mem_en_ctx2;
wire [5:0] MEMC53_start_addr_ctx2;
wire [0:0] MEMC53_stride_ctx2;
wire [31:0] MEMC53_data_in_ctx1;
wire [31:0] MEMC53_data_in_ctx2;
wire [31:0] MEMC53_data_out_ctx1;
wire [31:0] MEMC53_data_out_ctx2;
wire [63:0] MEMC53_burst_count_ctx1;
wire [63:0] MEMC53_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC53(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC53_data_from_Core),
.data_to_Core(MEMC53_data_to_Core),
.valid_ctx1(MEMC53_valid_ctx1),
.addr_out_ctx1(MEMC53_addr_out_ctx1),
.write_en_ctx1(MEMC53_write_en_ctx1),
.start_addr_ctx1(MEMC53_start_addr_ctx1),
.stride_ctx1(MEMC53_stride_ctx1),
.burst_count_ctx1(MEMC53_burst_count_ctx1),
.valid_ctx2(MEMC53_valid_ctx2),
.addr_out_ctx2(MEMC53_addr_out_ctx2),
.write_en_ctx2(MEMC53_write_en_ctx2),
.start_addr_ctx2(MEMC53_start_addr_ctx2),
.stride_ctx2(MEMC53_stride_ctx2),
.burst_count_ctx2(MEMC53_burst_count_ctx2),
.data_in_ctx1(MEMC53_data_in_ctx1),
.data_in_ctx2(MEMC53_data_in_ctx2),
.data_out_ctx1(MEMC53_data_out_ctx1),
.data_out_ctx2(MEMC53_data_out_ctx2),
.write_mem_en_ctx1(MEMC53_write_mem_en_ctx1),
.mem_en_ctx1(MEMC53_mem_en_ctx1),.write_mem_en_ctx2(MEMC53_write_mem_en_ctx2),
.mem_en_ctx2(MEMC53_mem_en_ctx2));

defparam MEMC53.DATA_WIDTH = 32;
defparam MEMC53.ADDR_WIDTH = 6;
defparam MEMC53.STRIDE_WIDTH = 1;
wire MEMC54_valid_ctx1;
wire MEMC54_valid_ctx2;
wire [31:0] MEMC54_data_from_Core;
wire [31:0] MEMC54_data_to_Core;
wire [5:0] MEMC54_addr_out_ctx1;
wire MEMC54_write_en_ctx1;
wire MEMC54_write_mem_en_ctx1;
wire MEMC54_mem_en_ctx1;
wire [5:0] MEMC54_start_addr_ctx1;
wire [0:0] MEMC54_stride_ctx1;
wire [5:0] MEMC54_addr_out_ctx2;
wire MEMC54_write_en_ctx2;
wire MEMC54_write_mem_en_ctx2;
wire MEMC54_mem_en_ctx2;
wire [5:0] MEMC54_start_addr_ctx2;
wire [0:0] MEMC54_stride_ctx2;
wire [31:0] MEMC54_data_in_ctx1;
wire [31:0] MEMC54_data_in_ctx2;
wire [31:0] MEMC54_data_out_ctx1;
wire [31:0] MEMC54_data_out_ctx2;
wire [63:0] MEMC54_burst_count_ctx1;
wire [63:0] MEMC54_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC54(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC54_data_from_Core),
.data_to_Core(MEMC54_data_to_Core),
.valid_ctx1(MEMC54_valid_ctx1),
.addr_out_ctx1(MEMC54_addr_out_ctx1),
.write_en_ctx1(MEMC54_write_en_ctx1),
.start_addr_ctx1(MEMC54_start_addr_ctx1),
.stride_ctx1(MEMC54_stride_ctx1),
.burst_count_ctx1(MEMC54_burst_count_ctx1),
.valid_ctx2(MEMC54_valid_ctx2),
.addr_out_ctx2(MEMC54_addr_out_ctx2),
.write_en_ctx2(MEMC54_write_en_ctx2),
.start_addr_ctx2(MEMC54_start_addr_ctx2),
.stride_ctx2(MEMC54_stride_ctx2),
.burst_count_ctx2(MEMC54_burst_count_ctx2),
.data_in_ctx1(MEMC54_data_in_ctx1),
.data_in_ctx2(MEMC54_data_in_ctx2),
.data_out_ctx1(MEMC54_data_out_ctx1),
.data_out_ctx2(MEMC54_data_out_ctx2),
.write_mem_en_ctx1(MEMC54_write_mem_en_ctx1),
.mem_en_ctx1(MEMC54_mem_en_ctx1),.write_mem_en_ctx2(MEMC54_write_mem_en_ctx2),
.mem_en_ctx2(MEMC54_mem_en_ctx2));

defparam MEMC54.DATA_WIDTH = 32;
defparam MEMC54.ADDR_WIDTH = 6;
defparam MEMC54.STRIDE_WIDTH = 1;
wire MEMC55_valid_ctx1;
wire MEMC55_valid_ctx2;
wire [31:0] MEMC55_data_from_Core;
wire [31:0] MEMC55_data_to_Core;
wire [5:0] MEMC55_addr_out_ctx1;
wire MEMC55_write_en_ctx1;
wire MEMC55_write_mem_en_ctx1;
wire MEMC55_mem_en_ctx1;
wire [5:0] MEMC55_start_addr_ctx1;
wire [0:0] MEMC55_stride_ctx1;
wire [5:0] MEMC55_addr_out_ctx2;
wire MEMC55_write_en_ctx2;
wire MEMC55_write_mem_en_ctx2;
wire MEMC55_mem_en_ctx2;
wire [5:0] MEMC55_start_addr_ctx2;
wire [0:0] MEMC55_stride_ctx2;
wire [31:0] MEMC55_data_in_ctx1;
wire [31:0] MEMC55_data_in_ctx2;
wire [31:0] MEMC55_data_out_ctx1;
wire [31:0] MEMC55_data_out_ctx2;
wire [63:0] MEMC55_burst_count_ctx1;
wire [63:0] MEMC55_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC55(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC55_data_from_Core),
.data_to_Core(MEMC55_data_to_Core),
.valid_ctx1(MEMC55_valid_ctx1),
.addr_out_ctx1(MEMC55_addr_out_ctx1),
.write_en_ctx1(MEMC55_write_en_ctx1),
.start_addr_ctx1(MEMC55_start_addr_ctx1),
.stride_ctx1(MEMC55_stride_ctx1),
.burst_count_ctx1(MEMC55_burst_count_ctx1),
.valid_ctx2(MEMC55_valid_ctx2),
.addr_out_ctx2(MEMC55_addr_out_ctx2),
.write_en_ctx2(MEMC55_write_en_ctx2),
.start_addr_ctx2(MEMC55_start_addr_ctx2),
.stride_ctx2(MEMC55_stride_ctx2),
.burst_count_ctx2(MEMC55_burst_count_ctx2),
.data_in_ctx1(MEMC55_data_in_ctx1),
.data_in_ctx2(MEMC55_data_in_ctx2),
.data_out_ctx1(MEMC55_data_out_ctx1),
.data_out_ctx2(MEMC55_data_out_ctx2),
.write_mem_en_ctx1(MEMC55_write_mem_en_ctx1),
.mem_en_ctx1(MEMC55_mem_en_ctx1),.write_mem_en_ctx2(MEMC55_write_mem_en_ctx2),
.mem_en_ctx2(MEMC55_mem_en_ctx2));

defparam MEMC55.DATA_WIDTH = 32;
defparam MEMC55.ADDR_WIDTH = 6;
defparam MEMC55.STRIDE_WIDTH = 1;
wire MEMC56_valid_ctx1;
wire MEMC56_valid_ctx2;
wire [31:0] MEMC56_data_from_Core;
wire [31:0] MEMC56_data_to_Core;
wire [5:0] MEMC56_addr_out_ctx1;
wire MEMC56_write_en_ctx1;
wire MEMC56_write_mem_en_ctx1;
wire MEMC56_mem_en_ctx1;
wire [5:0] MEMC56_start_addr_ctx1;
wire [0:0] MEMC56_stride_ctx1;
wire [5:0] MEMC56_addr_out_ctx2;
wire MEMC56_write_en_ctx2;
wire MEMC56_write_mem_en_ctx2;
wire MEMC56_mem_en_ctx2;
wire [5:0] MEMC56_start_addr_ctx2;
wire [0:0] MEMC56_stride_ctx2;
wire [31:0] MEMC56_data_in_ctx1;
wire [31:0] MEMC56_data_in_ctx2;
wire [31:0] MEMC56_data_out_ctx1;
wire [31:0] MEMC56_data_out_ctx2;
wire [63:0] MEMC56_burst_count_ctx1;
wire [63:0] MEMC56_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC56(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC56_data_from_Core),
.data_to_Core(MEMC56_data_to_Core),
.valid_ctx1(MEMC56_valid_ctx1),
.addr_out_ctx1(MEMC56_addr_out_ctx1),
.write_en_ctx1(MEMC56_write_en_ctx1),
.start_addr_ctx1(MEMC56_start_addr_ctx1),
.stride_ctx1(MEMC56_stride_ctx1),
.burst_count_ctx1(MEMC56_burst_count_ctx1),
.valid_ctx2(MEMC56_valid_ctx2),
.addr_out_ctx2(MEMC56_addr_out_ctx2),
.write_en_ctx2(MEMC56_write_en_ctx2),
.start_addr_ctx2(MEMC56_start_addr_ctx2),
.stride_ctx2(MEMC56_stride_ctx2),
.burst_count_ctx2(MEMC56_burst_count_ctx2),
.data_in_ctx1(MEMC56_data_in_ctx1),
.data_in_ctx2(MEMC56_data_in_ctx2),
.data_out_ctx1(MEMC56_data_out_ctx1),
.data_out_ctx2(MEMC56_data_out_ctx2),
.write_mem_en_ctx1(MEMC56_write_mem_en_ctx1),
.mem_en_ctx1(MEMC56_mem_en_ctx1),.write_mem_en_ctx2(MEMC56_write_mem_en_ctx2),
.mem_en_ctx2(MEMC56_mem_en_ctx2));

defparam MEMC56.DATA_WIDTH = 32;
defparam MEMC56.ADDR_WIDTH = 6;
defparam MEMC56.STRIDE_WIDTH = 1;
wire MEMC57_valid_ctx1;
wire MEMC57_valid_ctx2;
wire [31:0] MEMC57_data_from_Core;
wire [31:0] MEMC57_data_to_Core;
wire [5:0] MEMC57_addr_out_ctx1;
wire MEMC57_write_en_ctx1;
wire MEMC57_write_mem_en_ctx1;
wire MEMC57_mem_en_ctx1;
wire [5:0] MEMC57_start_addr_ctx1;
wire [0:0] MEMC57_stride_ctx1;
wire [5:0] MEMC57_addr_out_ctx2;
wire MEMC57_write_en_ctx2;
wire MEMC57_write_mem_en_ctx2;
wire MEMC57_mem_en_ctx2;
wire [5:0] MEMC57_start_addr_ctx2;
wire [0:0] MEMC57_stride_ctx2;
wire [31:0] MEMC57_data_in_ctx1;
wire [31:0] MEMC57_data_in_ctx2;
wire [31:0] MEMC57_data_out_ctx1;
wire [31:0] MEMC57_data_out_ctx2;
wire [63:0] MEMC57_burst_count_ctx1;
wire [63:0] MEMC57_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC57(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC57_data_from_Core),
.data_to_Core(MEMC57_data_to_Core),
.valid_ctx1(MEMC57_valid_ctx1),
.addr_out_ctx1(MEMC57_addr_out_ctx1),
.write_en_ctx1(MEMC57_write_en_ctx1),
.start_addr_ctx1(MEMC57_start_addr_ctx1),
.stride_ctx1(MEMC57_stride_ctx1),
.burst_count_ctx1(MEMC57_burst_count_ctx1),
.valid_ctx2(MEMC57_valid_ctx2),
.addr_out_ctx2(MEMC57_addr_out_ctx2),
.write_en_ctx2(MEMC57_write_en_ctx2),
.start_addr_ctx2(MEMC57_start_addr_ctx2),
.stride_ctx2(MEMC57_stride_ctx2),
.burst_count_ctx2(MEMC57_burst_count_ctx2),
.data_in_ctx1(MEMC57_data_in_ctx1),
.data_in_ctx2(MEMC57_data_in_ctx2),
.data_out_ctx1(MEMC57_data_out_ctx1),
.data_out_ctx2(MEMC57_data_out_ctx2),
.write_mem_en_ctx1(MEMC57_write_mem_en_ctx1),
.mem_en_ctx1(MEMC57_mem_en_ctx1),.write_mem_en_ctx2(MEMC57_write_mem_en_ctx2),
.mem_en_ctx2(MEMC57_mem_en_ctx2));

defparam MEMC57.DATA_WIDTH = 32;
defparam MEMC57.ADDR_WIDTH = 6;
defparam MEMC57.STRIDE_WIDTH = 1;
wire MEMC58_valid_ctx1;
wire MEMC58_valid_ctx2;
wire [31:0] MEMC58_data_from_Core;
wire [31:0] MEMC58_data_to_Core;
wire [5:0] MEMC58_addr_out_ctx1;
wire MEMC58_write_en_ctx1;
wire MEMC58_write_mem_en_ctx1;
wire MEMC58_mem_en_ctx1;
wire [5:0] MEMC58_start_addr_ctx1;
wire [0:0] MEMC58_stride_ctx1;
wire [5:0] MEMC58_addr_out_ctx2;
wire MEMC58_write_en_ctx2;
wire MEMC58_write_mem_en_ctx2;
wire MEMC58_mem_en_ctx2;
wire [5:0] MEMC58_start_addr_ctx2;
wire [0:0] MEMC58_stride_ctx2;
wire [31:0] MEMC58_data_in_ctx1;
wire [31:0] MEMC58_data_in_ctx2;
wire [31:0] MEMC58_data_out_ctx1;
wire [31:0] MEMC58_data_out_ctx2;
wire [63:0] MEMC58_burst_count_ctx1;
wire [63:0] MEMC58_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC58(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC58_data_from_Core),
.data_to_Core(MEMC58_data_to_Core),
.valid_ctx1(MEMC58_valid_ctx1),
.addr_out_ctx1(MEMC58_addr_out_ctx1),
.write_en_ctx1(MEMC58_write_en_ctx1),
.start_addr_ctx1(MEMC58_start_addr_ctx1),
.stride_ctx1(MEMC58_stride_ctx1),
.burst_count_ctx1(MEMC58_burst_count_ctx1),
.valid_ctx2(MEMC58_valid_ctx2),
.addr_out_ctx2(MEMC58_addr_out_ctx2),
.write_en_ctx2(MEMC58_write_en_ctx2),
.start_addr_ctx2(MEMC58_start_addr_ctx2),
.stride_ctx2(MEMC58_stride_ctx2),
.burst_count_ctx2(MEMC58_burst_count_ctx2),
.data_in_ctx1(MEMC58_data_in_ctx1),
.data_in_ctx2(MEMC58_data_in_ctx2),
.data_out_ctx1(MEMC58_data_out_ctx1),
.data_out_ctx2(MEMC58_data_out_ctx2),
.write_mem_en_ctx1(MEMC58_write_mem_en_ctx1),
.mem_en_ctx1(MEMC58_mem_en_ctx1),.write_mem_en_ctx2(MEMC58_write_mem_en_ctx2),
.mem_en_ctx2(MEMC58_mem_en_ctx2));

defparam MEMC58.DATA_WIDTH = 32;
defparam MEMC58.ADDR_WIDTH = 6;
defparam MEMC58.STRIDE_WIDTH = 1;
wire MEMC59_valid_ctx1;
wire MEMC59_valid_ctx2;
wire [31:0] MEMC59_data_from_Core;
wire [31:0] MEMC59_data_to_Core;
wire [5:0] MEMC59_addr_out_ctx1;
wire MEMC59_write_en_ctx1;
wire MEMC59_write_mem_en_ctx1;
wire MEMC59_mem_en_ctx1;
wire [5:0] MEMC59_start_addr_ctx1;
wire [0:0] MEMC59_stride_ctx1;
wire [5:0] MEMC59_addr_out_ctx2;
wire MEMC59_write_en_ctx2;
wire MEMC59_write_mem_en_ctx2;
wire MEMC59_mem_en_ctx2;
wire [5:0] MEMC59_start_addr_ctx2;
wire [0:0] MEMC59_stride_ctx2;
wire [31:0] MEMC59_data_in_ctx1;
wire [31:0] MEMC59_data_in_ctx2;
wire [31:0] MEMC59_data_out_ctx1;
wire [31:0] MEMC59_data_out_ctx2;
wire [63:0] MEMC59_burst_count_ctx1;
wire [63:0] MEMC59_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC59(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC59_data_from_Core),
.data_to_Core(MEMC59_data_to_Core),
.valid_ctx1(MEMC59_valid_ctx1),
.addr_out_ctx1(MEMC59_addr_out_ctx1),
.write_en_ctx1(MEMC59_write_en_ctx1),
.start_addr_ctx1(MEMC59_start_addr_ctx1),
.stride_ctx1(MEMC59_stride_ctx1),
.burst_count_ctx1(MEMC59_burst_count_ctx1),
.valid_ctx2(MEMC59_valid_ctx2),
.addr_out_ctx2(MEMC59_addr_out_ctx2),
.write_en_ctx2(MEMC59_write_en_ctx2),
.start_addr_ctx2(MEMC59_start_addr_ctx2),
.stride_ctx2(MEMC59_stride_ctx2),
.burst_count_ctx2(MEMC59_burst_count_ctx2),
.data_in_ctx1(MEMC59_data_in_ctx1),
.data_in_ctx2(MEMC59_data_in_ctx2),
.data_out_ctx1(MEMC59_data_out_ctx1),
.data_out_ctx2(MEMC59_data_out_ctx2),
.write_mem_en_ctx1(MEMC59_write_mem_en_ctx1),
.mem_en_ctx1(MEMC59_mem_en_ctx1),.write_mem_en_ctx2(MEMC59_write_mem_en_ctx2),
.mem_en_ctx2(MEMC59_mem_en_ctx2));

defparam MEMC59.DATA_WIDTH = 32;
defparam MEMC59.ADDR_WIDTH = 6;
defparam MEMC59.STRIDE_WIDTH = 1;
wire MEMC60_valid_ctx1;
wire MEMC60_valid_ctx2;
wire [31:0] MEMC60_data_from_Core;
wire [31:0] MEMC60_data_to_Core;
wire [5:0] MEMC60_addr_out_ctx1;
wire MEMC60_write_en_ctx1;
wire MEMC60_write_mem_en_ctx1;
wire MEMC60_mem_en_ctx1;
wire [5:0] MEMC60_start_addr_ctx1;
wire [0:0] MEMC60_stride_ctx1;
wire [5:0] MEMC60_addr_out_ctx2;
wire MEMC60_write_en_ctx2;
wire MEMC60_write_mem_en_ctx2;
wire MEMC60_mem_en_ctx2;
wire [5:0] MEMC60_start_addr_ctx2;
wire [0:0] MEMC60_stride_ctx2;
wire [31:0] MEMC60_data_in_ctx1;
wire [31:0] MEMC60_data_in_ctx2;
wire [31:0] MEMC60_data_out_ctx1;
wire [31:0] MEMC60_data_out_ctx2;
wire [63:0] MEMC60_burst_count_ctx1;
wire [63:0] MEMC60_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC60(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC60_data_from_Core),
.data_to_Core(MEMC60_data_to_Core),
.valid_ctx1(MEMC60_valid_ctx1),
.addr_out_ctx1(MEMC60_addr_out_ctx1),
.write_en_ctx1(MEMC60_write_en_ctx1),
.start_addr_ctx1(MEMC60_start_addr_ctx1),
.stride_ctx1(MEMC60_stride_ctx1),
.burst_count_ctx1(MEMC60_burst_count_ctx1),
.valid_ctx2(MEMC60_valid_ctx2),
.addr_out_ctx2(MEMC60_addr_out_ctx2),
.write_en_ctx2(MEMC60_write_en_ctx2),
.start_addr_ctx2(MEMC60_start_addr_ctx2),
.stride_ctx2(MEMC60_stride_ctx2),
.burst_count_ctx2(MEMC60_burst_count_ctx2),
.data_in_ctx1(MEMC60_data_in_ctx1),
.data_in_ctx2(MEMC60_data_in_ctx2),
.data_out_ctx1(MEMC60_data_out_ctx1),
.data_out_ctx2(MEMC60_data_out_ctx2),
.write_mem_en_ctx1(MEMC60_write_mem_en_ctx1),
.mem_en_ctx1(MEMC60_mem_en_ctx1),.write_mem_en_ctx2(MEMC60_write_mem_en_ctx2),
.mem_en_ctx2(MEMC60_mem_en_ctx2));

defparam MEMC60.DATA_WIDTH = 32;
defparam MEMC60.ADDR_WIDTH = 6;
defparam MEMC60.STRIDE_WIDTH = 1;
wire MEMC61_valid_ctx1;
wire MEMC61_valid_ctx2;
wire [31:0] MEMC61_data_from_Core;
wire [31:0] MEMC61_data_to_Core;
wire [5:0] MEMC61_addr_out_ctx1;
wire MEMC61_write_en_ctx1;
wire MEMC61_write_mem_en_ctx1;
wire MEMC61_mem_en_ctx1;
wire [5:0] MEMC61_start_addr_ctx1;
wire [0:0] MEMC61_stride_ctx1;
wire [5:0] MEMC61_addr_out_ctx2;
wire MEMC61_write_en_ctx2;
wire MEMC61_write_mem_en_ctx2;
wire MEMC61_mem_en_ctx2;
wire [5:0] MEMC61_start_addr_ctx2;
wire [0:0] MEMC61_stride_ctx2;
wire [31:0] MEMC61_data_in_ctx1;
wire [31:0] MEMC61_data_in_ctx2;
wire [31:0] MEMC61_data_out_ctx1;
wire [31:0] MEMC61_data_out_ctx2;
wire [63:0] MEMC61_burst_count_ctx1;
wire [63:0] MEMC61_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC61(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC61_data_from_Core),
.data_to_Core(MEMC61_data_to_Core),
.valid_ctx1(MEMC61_valid_ctx1),
.addr_out_ctx1(MEMC61_addr_out_ctx1),
.write_en_ctx1(MEMC61_write_en_ctx1),
.start_addr_ctx1(MEMC61_start_addr_ctx1),
.stride_ctx1(MEMC61_stride_ctx1),
.burst_count_ctx1(MEMC61_burst_count_ctx1),
.valid_ctx2(MEMC61_valid_ctx2),
.addr_out_ctx2(MEMC61_addr_out_ctx2),
.write_en_ctx2(MEMC61_write_en_ctx2),
.start_addr_ctx2(MEMC61_start_addr_ctx2),
.stride_ctx2(MEMC61_stride_ctx2),
.burst_count_ctx2(MEMC61_burst_count_ctx2),
.data_in_ctx1(MEMC61_data_in_ctx1),
.data_in_ctx2(MEMC61_data_in_ctx2),
.data_out_ctx1(MEMC61_data_out_ctx1),
.data_out_ctx2(MEMC61_data_out_ctx2),
.write_mem_en_ctx1(MEMC61_write_mem_en_ctx1),
.mem_en_ctx1(MEMC61_mem_en_ctx1),.write_mem_en_ctx2(MEMC61_write_mem_en_ctx2),
.mem_en_ctx2(MEMC61_mem_en_ctx2));

defparam MEMC61.DATA_WIDTH = 32;
defparam MEMC61.ADDR_WIDTH = 6;
defparam MEMC61.STRIDE_WIDTH = 1;
wire MEMC62_valid_ctx1;
wire MEMC62_valid_ctx2;
wire [31:0] MEMC62_data_from_Core;
wire [31:0] MEMC62_data_to_Core;
wire [5:0] MEMC62_addr_out_ctx1;
wire MEMC62_write_en_ctx1;
wire MEMC62_write_mem_en_ctx1;
wire MEMC62_mem_en_ctx1;
wire [5:0] MEMC62_start_addr_ctx1;
wire [0:0] MEMC62_stride_ctx1;
wire [5:0] MEMC62_addr_out_ctx2;
wire MEMC62_write_en_ctx2;
wire MEMC62_write_mem_en_ctx2;
wire MEMC62_mem_en_ctx2;
wire [5:0] MEMC62_start_addr_ctx2;
wire [0:0] MEMC62_stride_ctx2;
wire [31:0] MEMC62_data_in_ctx1;
wire [31:0] MEMC62_data_in_ctx2;
wire [31:0] MEMC62_data_out_ctx1;
wire [31:0] MEMC62_data_out_ctx2;
wire [63:0] MEMC62_burst_count_ctx1;
wire [63:0] MEMC62_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC62(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC62_data_from_Core),
.data_to_Core(MEMC62_data_to_Core),
.valid_ctx1(MEMC62_valid_ctx1),
.addr_out_ctx1(MEMC62_addr_out_ctx1),
.write_en_ctx1(MEMC62_write_en_ctx1),
.start_addr_ctx1(MEMC62_start_addr_ctx1),
.stride_ctx1(MEMC62_stride_ctx1),
.burst_count_ctx1(MEMC62_burst_count_ctx1),
.valid_ctx2(MEMC62_valid_ctx2),
.addr_out_ctx2(MEMC62_addr_out_ctx2),
.write_en_ctx2(MEMC62_write_en_ctx2),
.start_addr_ctx2(MEMC62_start_addr_ctx2),
.stride_ctx2(MEMC62_stride_ctx2),
.burst_count_ctx2(MEMC62_burst_count_ctx2),
.data_in_ctx1(MEMC62_data_in_ctx1),
.data_in_ctx2(MEMC62_data_in_ctx2),
.data_out_ctx1(MEMC62_data_out_ctx1),
.data_out_ctx2(MEMC62_data_out_ctx2),
.write_mem_en_ctx1(MEMC62_write_mem_en_ctx1),
.mem_en_ctx1(MEMC62_mem_en_ctx1),.write_mem_en_ctx2(MEMC62_write_mem_en_ctx2),
.mem_en_ctx2(MEMC62_mem_en_ctx2));

defparam MEMC62.DATA_WIDTH = 32;
defparam MEMC62.ADDR_WIDTH = 6;
defparam MEMC62.STRIDE_WIDTH = 1;
wire MEMC63_valid_ctx1;
wire MEMC63_valid_ctx2;
wire [31:0] MEMC63_data_from_Core;
wire [31:0] MEMC63_data_to_Core;
wire [5:0] MEMC63_addr_out_ctx1;
wire MEMC63_write_en_ctx1;
wire MEMC63_write_mem_en_ctx1;
wire MEMC63_mem_en_ctx1;
wire [5:0] MEMC63_start_addr_ctx1;
wire [0:0] MEMC63_stride_ctx1;
wire [5:0] MEMC63_addr_out_ctx2;
wire MEMC63_write_en_ctx2;
wire MEMC63_write_mem_en_ctx2;
wire MEMC63_mem_en_ctx2;
wire [5:0] MEMC63_start_addr_ctx2;
wire [0:0] MEMC63_stride_ctx2;
wire [31:0] MEMC63_data_in_ctx1;
wire [31:0] MEMC63_data_in_ctx2;
wire [31:0] MEMC63_data_out_ctx1;
wire [31:0] MEMC63_data_out_ctx2;
wire [63:0] MEMC63_burst_count_ctx1;
wire [63:0] MEMC63_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC63(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC63_data_from_Core),
.data_to_Core(MEMC63_data_to_Core),
.valid_ctx1(MEMC63_valid_ctx1),
.addr_out_ctx1(MEMC63_addr_out_ctx1),
.write_en_ctx1(MEMC63_write_en_ctx1),
.start_addr_ctx1(MEMC63_start_addr_ctx1),
.stride_ctx1(MEMC63_stride_ctx1),
.burst_count_ctx1(MEMC63_burst_count_ctx1),
.valid_ctx2(MEMC63_valid_ctx2),
.addr_out_ctx2(MEMC63_addr_out_ctx2),
.write_en_ctx2(MEMC63_write_en_ctx2),
.start_addr_ctx2(MEMC63_start_addr_ctx2),
.stride_ctx2(MEMC63_stride_ctx2),
.burst_count_ctx2(MEMC63_burst_count_ctx2),
.data_in_ctx1(MEMC63_data_in_ctx1),
.data_in_ctx2(MEMC63_data_in_ctx2),
.data_out_ctx1(MEMC63_data_out_ctx1),
.data_out_ctx2(MEMC63_data_out_ctx2),
.write_mem_en_ctx1(MEMC63_write_mem_en_ctx1),
.mem_en_ctx1(MEMC63_mem_en_ctx1),.write_mem_en_ctx2(MEMC63_write_mem_en_ctx2),
.mem_en_ctx2(MEMC63_mem_en_ctx2));

defparam MEMC63.DATA_WIDTH = 32;
defparam MEMC63.ADDR_WIDTH = 6;
defparam MEMC63.STRIDE_WIDTH = 1;
wire MEMC64_valid_ctx1;
wire MEMC64_valid_ctx2;
wire [31:0] MEMC64_data_from_Core;
wire [31:0] MEMC64_data_to_Core;
wire [5:0] MEMC64_addr_out_ctx1;
wire MEMC64_write_en_ctx1;
wire MEMC64_write_mem_en_ctx1;
wire MEMC64_mem_en_ctx1;
wire [5:0] MEMC64_start_addr_ctx1;
wire [0:0] MEMC64_stride_ctx1;
wire [5:0] MEMC64_addr_out_ctx2;
wire MEMC64_write_en_ctx2;
wire MEMC64_write_mem_en_ctx2;
wire MEMC64_mem_en_ctx2;
wire [5:0] MEMC64_start_addr_ctx2;
wire [0:0] MEMC64_stride_ctx2;
wire [31:0] MEMC64_data_in_ctx1;
wire [31:0] MEMC64_data_in_ctx2;
wire [31:0] MEMC64_data_out_ctx1;
wire [31:0] MEMC64_data_out_ctx2;
wire [63:0] MEMC64_burst_count_ctx1;
wire [63:0] MEMC64_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC64(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC64_data_from_Core),
.data_to_Core(MEMC64_data_to_Core),
.valid_ctx1(MEMC64_valid_ctx1),
.addr_out_ctx1(MEMC64_addr_out_ctx1),
.write_en_ctx1(MEMC64_write_en_ctx1),
.start_addr_ctx1(MEMC64_start_addr_ctx1),
.stride_ctx1(MEMC64_stride_ctx1),
.burst_count_ctx1(MEMC64_burst_count_ctx1),
.valid_ctx2(MEMC64_valid_ctx2),
.addr_out_ctx2(MEMC64_addr_out_ctx2),
.write_en_ctx2(MEMC64_write_en_ctx2),
.start_addr_ctx2(MEMC64_start_addr_ctx2),
.stride_ctx2(MEMC64_stride_ctx2),
.burst_count_ctx2(MEMC64_burst_count_ctx2),
.data_in_ctx1(MEMC64_data_in_ctx1),
.data_in_ctx2(MEMC64_data_in_ctx2),
.data_out_ctx1(MEMC64_data_out_ctx1),
.data_out_ctx2(MEMC64_data_out_ctx2),
.write_mem_en_ctx1(MEMC64_write_mem_en_ctx1),
.mem_en_ctx1(MEMC64_mem_en_ctx1),.write_mem_en_ctx2(MEMC64_write_mem_en_ctx2),
.mem_en_ctx2(MEMC64_mem_en_ctx2));

defparam MEMC64.DATA_WIDTH = 32;
defparam MEMC64.ADDR_WIDTH = 6;
defparam MEMC64.STRIDE_WIDTH = 1;
wire MEMC65_valid_ctx1;
wire MEMC65_valid_ctx2;
wire [31:0] MEMC65_data_from_Core;
wire [31:0] MEMC65_data_to_Core;
wire [5:0] MEMC65_addr_out_ctx1;
wire MEMC65_write_en_ctx1;
wire MEMC65_write_mem_en_ctx1;
wire MEMC65_mem_en_ctx1;
wire [5:0] MEMC65_start_addr_ctx1;
wire [0:0] MEMC65_stride_ctx1;
wire [5:0] MEMC65_addr_out_ctx2;
wire MEMC65_write_en_ctx2;
wire MEMC65_write_mem_en_ctx2;
wire MEMC65_mem_en_ctx2;
wire [5:0] MEMC65_start_addr_ctx2;
wire [0:0] MEMC65_stride_ctx2;
wire [31:0] MEMC65_data_in_ctx1;
wire [31:0] MEMC65_data_in_ctx2;
wire [31:0] MEMC65_data_out_ctx1;
wire [31:0] MEMC65_data_out_ctx2;
wire [63:0] MEMC65_burst_count_ctx1;
wire [63:0] MEMC65_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC65(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC65_data_from_Core),
.data_to_Core(MEMC65_data_to_Core),
.valid_ctx1(MEMC65_valid_ctx1),
.addr_out_ctx1(MEMC65_addr_out_ctx1),
.write_en_ctx1(MEMC65_write_en_ctx1),
.start_addr_ctx1(MEMC65_start_addr_ctx1),
.stride_ctx1(MEMC65_stride_ctx1),
.burst_count_ctx1(MEMC65_burst_count_ctx1),
.valid_ctx2(MEMC65_valid_ctx2),
.addr_out_ctx2(MEMC65_addr_out_ctx2),
.write_en_ctx2(MEMC65_write_en_ctx2),
.start_addr_ctx2(MEMC65_start_addr_ctx2),
.stride_ctx2(MEMC65_stride_ctx2),
.burst_count_ctx2(MEMC65_burst_count_ctx2),
.data_in_ctx1(MEMC65_data_in_ctx1),
.data_in_ctx2(MEMC65_data_in_ctx2),
.data_out_ctx1(MEMC65_data_out_ctx1),
.data_out_ctx2(MEMC65_data_out_ctx2),
.write_mem_en_ctx1(MEMC65_write_mem_en_ctx1),
.mem_en_ctx1(MEMC65_mem_en_ctx1),.write_mem_en_ctx2(MEMC65_write_mem_en_ctx2),
.mem_en_ctx2(MEMC65_mem_en_ctx2));

defparam MEMC65.DATA_WIDTH = 32;
defparam MEMC65.ADDR_WIDTH = 6;
defparam MEMC65.STRIDE_WIDTH = 1;
wire MEMC66_valid_ctx1;
wire MEMC66_valid_ctx2;
wire [31:0] MEMC66_data_from_Core;
wire [31:0] MEMC66_data_to_Core;
wire [5:0] MEMC66_addr_out_ctx1;
wire MEMC66_write_en_ctx1;
wire MEMC66_write_mem_en_ctx1;
wire MEMC66_mem_en_ctx1;
wire [5:0] MEMC66_start_addr_ctx1;
wire [0:0] MEMC66_stride_ctx1;
wire [5:0] MEMC66_addr_out_ctx2;
wire MEMC66_write_en_ctx2;
wire MEMC66_write_mem_en_ctx2;
wire MEMC66_mem_en_ctx2;
wire [5:0] MEMC66_start_addr_ctx2;
wire [0:0] MEMC66_stride_ctx2;
wire [31:0] MEMC66_data_in_ctx1;
wire [31:0] MEMC66_data_in_ctx2;
wire [31:0] MEMC66_data_out_ctx1;
wire [31:0] MEMC66_data_out_ctx2;
wire [63:0] MEMC66_burst_count_ctx1;
wire [63:0] MEMC66_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC66(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC66_data_from_Core),
.data_to_Core(MEMC66_data_to_Core),
.valid_ctx1(MEMC66_valid_ctx1),
.addr_out_ctx1(MEMC66_addr_out_ctx1),
.write_en_ctx1(MEMC66_write_en_ctx1),
.start_addr_ctx1(MEMC66_start_addr_ctx1),
.stride_ctx1(MEMC66_stride_ctx1),
.burst_count_ctx1(MEMC66_burst_count_ctx1),
.valid_ctx2(MEMC66_valid_ctx2),
.addr_out_ctx2(MEMC66_addr_out_ctx2),
.write_en_ctx2(MEMC66_write_en_ctx2),
.start_addr_ctx2(MEMC66_start_addr_ctx2),
.stride_ctx2(MEMC66_stride_ctx2),
.burst_count_ctx2(MEMC66_burst_count_ctx2),
.data_in_ctx1(MEMC66_data_in_ctx1),
.data_in_ctx2(MEMC66_data_in_ctx2),
.data_out_ctx1(MEMC66_data_out_ctx1),
.data_out_ctx2(MEMC66_data_out_ctx2),
.write_mem_en_ctx1(MEMC66_write_mem_en_ctx1),
.mem_en_ctx1(MEMC66_mem_en_ctx1),.write_mem_en_ctx2(MEMC66_write_mem_en_ctx2),
.mem_en_ctx2(MEMC66_mem_en_ctx2));

defparam MEMC66.DATA_WIDTH = 32;
defparam MEMC66.ADDR_WIDTH = 6;
defparam MEMC66.STRIDE_WIDTH = 1;
wire MEMC67_valid_ctx1;
wire MEMC67_valid_ctx2;
wire [31:0] MEMC67_data_from_Core;
wire [31:0] MEMC67_data_to_Core;
wire [5:0] MEMC67_addr_out_ctx1;
wire MEMC67_write_en_ctx1;
wire MEMC67_write_mem_en_ctx1;
wire MEMC67_mem_en_ctx1;
wire [5:0] MEMC67_start_addr_ctx1;
wire [0:0] MEMC67_stride_ctx1;
wire [5:0] MEMC67_addr_out_ctx2;
wire MEMC67_write_en_ctx2;
wire MEMC67_write_mem_en_ctx2;
wire MEMC67_mem_en_ctx2;
wire [5:0] MEMC67_start_addr_ctx2;
wire [0:0] MEMC67_stride_ctx2;
wire [31:0] MEMC67_data_in_ctx1;
wire [31:0] MEMC67_data_in_ctx2;
wire [31:0] MEMC67_data_out_ctx1;
wire [31:0] MEMC67_data_out_ctx2;
wire [63:0] MEMC67_burst_count_ctx1;
wire [63:0] MEMC67_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC67(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC67_data_from_Core),
.data_to_Core(MEMC67_data_to_Core),
.valid_ctx1(MEMC67_valid_ctx1),
.addr_out_ctx1(MEMC67_addr_out_ctx1),
.write_en_ctx1(MEMC67_write_en_ctx1),
.start_addr_ctx1(MEMC67_start_addr_ctx1),
.stride_ctx1(MEMC67_stride_ctx1),
.burst_count_ctx1(MEMC67_burst_count_ctx1),
.valid_ctx2(MEMC67_valid_ctx2),
.addr_out_ctx2(MEMC67_addr_out_ctx2),
.write_en_ctx2(MEMC67_write_en_ctx2),
.start_addr_ctx2(MEMC67_start_addr_ctx2),
.stride_ctx2(MEMC67_stride_ctx2),
.burst_count_ctx2(MEMC67_burst_count_ctx2),
.data_in_ctx1(MEMC67_data_in_ctx1),
.data_in_ctx2(MEMC67_data_in_ctx2),
.data_out_ctx1(MEMC67_data_out_ctx1),
.data_out_ctx2(MEMC67_data_out_ctx2),
.write_mem_en_ctx1(MEMC67_write_mem_en_ctx1),
.mem_en_ctx1(MEMC67_mem_en_ctx1),.write_mem_en_ctx2(MEMC67_write_mem_en_ctx2),
.mem_en_ctx2(MEMC67_mem_en_ctx2));

defparam MEMC67.DATA_WIDTH = 32;
defparam MEMC67.ADDR_WIDTH = 6;
defparam MEMC67.STRIDE_WIDTH = 1;
wire MEMC68_valid_ctx1;
wire MEMC68_valid_ctx2;
wire [31:0] MEMC68_data_from_Core;
wire [31:0] MEMC68_data_to_Core;
wire [5:0] MEMC68_addr_out_ctx1;
wire MEMC68_write_en_ctx1;
wire MEMC68_write_mem_en_ctx1;
wire MEMC68_mem_en_ctx1;
wire [5:0] MEMC68_start_addr_ctx1;
wire [0:0] MEMC68_stride_ctx1;
wire [5:0] MEMC68_addr_out_ctx2;
wire MEMC68_write_en_ctx2;
wire MEMC68_write_mem_en_ctx2;
wire MEMC68_mem_en_ctx2;
wire [5:0] MEMC68_start_addr_ctx2;
wire [0:0] MEMC68_stride_ctx2;
wire [31:0] MEMC68_data_in_ctx1;
wire [31:0] MEMC68_data_in_ctx2;
wire [31:0] MEMC68_data_out_ctx1;
wire [31:0] MEMC68_data_out_ctx2;
wire [63:0] MEMC68_burst_count_ctx1;
wire [63:0] MEMC68_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC68(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC68_data_from_Core),
.data_to_Core(MEMC68_data_to_Core),
.valid_ctx1(MEMC68_valid_ctx1),
.addr_out_ctx1(MEMC68_addr_out_ctx1),
.write_en_ctx1(MEMC68_write_en_ctx1),
.start_addr_ctx1(MEMC68_start_addr_ctx1),
.stride_ctx1(MEMC68_stride_ctx1),
.burst_count_ctx1(MEMC68_burst_count_ctx1),
.valid_ctx2(MEMC68_valid_ctx2),
.addr_out_ctx2(MEMC68_addr_out_ctx2),
.write_en_ctx2(MEMC68_write_en_ctx2),
.start_addr_ctx2(MEMC68_start_addr_ctx2),
.stride_ctx2(MEMC68_stride_ctx2),
.burst_count_ctx2(MEMC68_burst_count_ctx2),
.data_in_ctx1(MEMC68_data_in_ctx1),
.data_in_ctx2(MEMC68_data_in_ctx2),
.data_out_ctx1(MEMC68_data_out_ctx1),
.data_out_ctx2(MEMC68_data_out_ctx2),
.write_mem_en_ctx1(MEMC68_write_mem_en_ctx1),
.mem_en_ctx1(MEMC68_mem_en_ctx1),.write_mem_en_ctx2(MEMC68_write_mem_en_ctx2),
.mem_en_ctx2(MEMC68_mem_en_ctx2));

defparam MEMC68.DATA_WIDTH = 32;
defparam MEMC68.ADDR_WIDTH = 6;
defparam MEMC68.STRIDE_WIDTH = 1;
wire MEMC69_valid_ctx1;
wire MEMC69_valid_ctx2;
wire [31:0] MEMC69_data_from_Core;
wire [31:0] MEMC69_data_to_Core;
wire [5:0] MEMC69_addr_out_ctx1;
wire MEMC69_write_en_ctx1;
wire MEMC69_write_mem_en_ctx1;
wire MEMC69_mem_en_ctx1;
wire [5:0] MEMC69_start_addr_ctx1;
wire [0:0] MEMC69_stride_ctx1;
wire [5:0] MEMC69_addr_out_ctx2;
wire MEMC69_write_en_ctx2;
wire MEMC69_write_mem_en_ctx2;
wire MEMC69_mem_en_ctx2;
wire [5:0] MEMC69_start_addr_ctx2;
wire [0:0] MEMC69_stride_ctx2;
wire [31:0] MEMC69_data_in_ctx1;
wire [31:0] MEMC69_data_in_ctx2;
wire [31:0] MEMC69_data_out_ctx1;
wire [31:0] MEMC69_data_out_ctx2;
wire [63:0] MEMC69_burst_count_ctx1;
wire [63:0] MEMC69_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC69(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC69_data_from_Core),
.data_to_Core(MEMC69_data_to_Core),
.valid_ctx1(MEMC69_valid_ctx1),
.addr_out_ctx1(MEMC69_addr_out_ctx1),
.write_en_ctx1(MEMC69_write_en_ctx1),
.start_addr_ctx1(MEMC69_start_addr_ctx1),
.stride_ctx1(MEMC69_stride_ctx1),
.burst_count_ctx1(MEMC69_burst_count_ctx1),
.valid_ctx2(MEMC69_valid_ctx2),
.addr_out_ctx2(MEMC69_addr_out_ctx2),
.write_en_ctx2(MEMC69_write_en_ctx2),
.start_addr_ctx2(MEMC69_start_addr_ctx2),
.stride_ctx2(MEMC69_stride_ctx2),
.burst_count_ctx2(MEMC69_burst_count_ctx2),
.data_in_ctx1(MEMC69_data_in_ctx1),
.data_in_ctx2(MEMC69_data_in_ctx2),
.data_out_ctx1(MEMC69_data_out_ctx1),
.data_out_ctx2(MEMC69_data_out_ctx2),
.write_mem_en_ctx1(MEMC69_write_mem_en_ctx1),
.mem_en_ctx1(MEMC69_mem_en_ctx1),.write_mem_en_ctx2(MEMC69_write_mem_en_ctx2),
.mem_en_ctx2(MEMC69_mem_en_ctx2));

defparam MEMC69.DATA_WIDTH = 32;
defparam MEMC69.ADDR_WIDTH = 6;
defparam MEMC69.STRIDE_WIDTH = 1;
wire MEMC70_valid_ctx1;
wire MEMC70_valid_ctx2;
wire [31:0] MEMC70_data_from_Core;
wire [31:0] MEMC70_data_to_Core;
wire [5:0] MEMC70_addr_out_ctx1;
wire MEMC70_write_en_ctx1;
wire MEMC70_write_mem_en_ctx1;
wire MEMC70_mem_en_ctx1;
wire [5:0] MEMC70_start_addr_ctx1;
wire [0:0] MEMC70_stride_ctx1;
wire [5:0] MEMC70_addr_out_ctx2;
wire MEMC70_write_en_ctx2;
wire MEMC70_write_mem_en_ctx2;
wire MEMC70_mem_en_ctx2;
wire [5:0] MEMC70_start_addr_ctx2;
wire [0:0] MEMC70_stride_ctx2;
wire [31:0] MEMC70_data_in_ctx1;
wire [31:0] MEMC70_data_in_ctx2;
wire [31:0] MEMC70_data_out_ctx1;
wire [31:0] MEMC70_data_out_ctx2;
wire [63:0] MEMC70_burst_count_ctx1;
wire [63:0] MEMC70_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC70(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC70_data_from_Core),
.data_to_Core(MEMC70_data_to_Core),
.valid_ctx1(MEMC70_valid_ctx1),
.addr_out_ctx1(MEMC70_addr_out_ctx1),
.write_en_ctx1(MEMC70_write_en_ctx1),
.start_addr_ctx1(MEMC70_start_addr_ctx1),
.stride_ctx1(MEMC70_stride_ctx1),
.burst_count_ctx1(MEMC70_burst_count_ctx1),
.valid_ctx2(MEMC70_valid_ctx2),
.addr_out_ctx2(MEMC70_addr_out_ctx2),
.write_en_ctx2(MEMC70_write_en_ctx2),
.start_addr_ctx2(MEMC70_start_addr_ctx2),
.stride_ctx2(MEMC70_stride_ctx2),
.burst_count_ctx2(MEMC70_burst_count_ctx2),
.data_in_ctx1(MEMC70_data_in_ctx1),
.data_in_ctx2(MEMC70_data_in_ctx2),
.data_out_ctx1(MEMC70_data_out_ctx1),
.data_out_ctx2(MEMC70_data_out_ctx2),
.write_mem_en_ctx1(MEMC70_write_mem_en_ctx1),
.mem_en_ctx1(MEMC70_mem_en_ctx1),.write_mem_en_ctx2(MEMC70_write_mem_en_ctx2),
.mem_en_ctx2(MEMC70_mem_en_ctx2));

defparam MEMC70.DATA_WIDTH = 32;
defparam MEMC70.ADDR_WIDTH = 6;
defparam MEMC70.STRIDE_WIDTH = 1;
wire MEMC71_valid_ctx1;
wire MEMC71_valid_ctx2;
wire [31:0] MEMC71_data_from_Core;
wire [31:0] MEMC71_data_to_Core;
wire [5:0] MEMC71_addr_out_ctx1;
wire MEMC71_write_en_ctx1;
wire MEMC71_write_mem_en_ctx1;
wire MEMC71_mem_en_ctx1;
wire [5:0] MEMC71_start_addr_ctx1;
wire [0:0] MEMC71_stride_ctx1;
wire [5:0] MEMC71_addr_out_ctx2;
wire MEMC71_write_en_ctx2;
wire MEMC71_write_mem_en_ctx2;
wire MEMC71_mem_en_ctx2;
wire [5:0] MEMC71_start_addr_ctx2;
wire [0:0] MEMC71_stride_ctx2;
wire [31:0] MEMC71_data_in_ctx1;
wire [31:0] MEMC71_data_in_ctx2;
wire [31:0] MEMC71_data_out_ctx1;
wire [31:0] MEMC71_data_out_ctx2;
wire [63:0] MEMC71_burst_count_ctx1;
wire [63:0] MEMC71_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC71(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC71_data_from_Core),
.data_to_Core(MEMC71_data_to_Core),
.valid_ctx1(MEMC71_valid_ctx1),
.addr_out_ctx1(MEMC71_addr_out_ctx1),
.write_en_ctx1(MEMC71_write_en_ctx1),
.start_addr_ctx1(MEMC71_start_addr_ctx1),
.stride_ctx1(MEMC71_stride_ctx1),
.burst_count_ctx1(MEMC71_burst_count_ctx1),
.valid_ctx2(MEMC71_valid_ctx2),
.addr_out_ctx2(MEMC71_addr_out_ctx2),
.write_en_ctx2(MEMC71_write_en_ctx2),
.start_addr_ctx2(MEMC71_start_addr_ctx2),
.stride_ctx2(MEMC71_stride_ctx2),
.burst_count_ctx2(MEMC71_burst_count_ctx2),
.data_in_ctx1(MEMC71_data_in_ctx1),
.data_in_ctx2(MEMC71_data_in_ctx2),
.data_out_ctx1(MEMC71_data_out_ctx1),
.data_out_ctx2(MEMC71_data_out_ctx2),
.write_mem_en_ctx1(MEMC71_write_mem_en_ctx1),
.mem_en_ctx1(MEMC71_mem_en_ctx1),.write_mem_en_ctx2(MEMC71_write_mem_en_ctx2),
.mem_en_ctx2(MEMC71_mem_en_ctx2));

defparam MEMC71.DATA_WIDTH = 32;
defparam MEMC71.ADDR_WIDTH = 6;
defparam MEMC71.STRIDE_WIDTH = 1;
wire MEMC72_valid_ctx1;
wire MEMC72_valid_ctx2;
wire [31:0] MEMC72_data_from_Core;
wire [31:0] MEMC72_data_to_Core;
wire [5:0] MEMC72_addr_out_ctx1;
wire MEMC72_write_en_ctx1;
wire MEMC72_write_mem_en_ctx1;
wire MEMC72_mem_en_ctx1;
wire [5:0] MEMC72_start_addr_ctx1;
wire [0:0] MEMC72_stride_ctx1;
wire [5:0] MEMC72_addr_out_ctx2;
wire MEMC72_write_en_ctx2;
wire MEMC72_write_mem_en_ctx2;
wire MEMC72_mem_en_ctx2;
wire [5:0] MEMC72_start_addr_ctx2;
wire [0:0] MEMC72_stride_ctx2;
wire [31:0] MEMC72_data_in_ctx1;
wire [31:0] MEMC72_data_in_ctx2;
wire [31:0] MEMC72_data_out_ctx1;
wire [31:0] MEMC72_data_out_ctx2;
wire [63:0] MEMC72_burst_count_ctx1;
wire [63:0] MEMC72_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC72(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC72_data_from_Core),
.data_to_Core(MEMC72_data_to_Core),
.valid_ctx1(MEMC72_valid_ctx1),
.addr_out_ctx1(MEMC72_addr_out_ctx1),
.write_en_ctx1(MEMC72_write_en_ctx1),
.start_addr_ctx1(MEMC72_start_addr_ctx1),
.stride_ctx1(MEMC72_stride_ctx1),
.burst_count_ctx1(MEMC72_burst_count_ctx1),
.valid_ctx2(MEMC72_valid_ctx2),
.addr_out_ctx2(MEMC72_addr_out_ctx2),
.write_en_ctx2(MEMC72_write_en_ctx2),
.start_addr_ctx2(MEMC72_start_addr_ctx2),
.stride_ctx2(MEMC72_stride_ctx2),
.burst_count_ctx2(MEMC72_burst_count_ctx2),
.data_in_ctx1(MEMC72_data_in_ctx1),
.data_in_ctx2(MEMC72_data_in_ctx2),
.data_out_ctx1(MEMC72_data_out_ctx1),
.data_out_ctx2(MEMC72_data_out_ctx2),
.write_mem_en_ctx1(MEMC72_write_mem_en_ctx1),
.mem_en_ctx1(MEMC72_mem_en_ctx1),.write_mem_en_ctx2(MEMC72_write_mem_en_ctx2),
.mem_en_ctx2(MEMC72_mem_en_ctx2));

defparam MEMC72.DATA_WIDTH = 32;
defparam MEMC72.ADDR_WIDTH = 6;
defparam MEMC72.STRIDE_WIDTH = 1;
wire MEMC73_valid_ctx1;
wire MEMC73_valid_ctx2;
wire [31:0] MEMC73_data_from_Core;
wire [31:0] MEMC73_data_to_Core;
wire [5:0] MEMC73_addr_out_ctx1;
wire MEMC73_write_en_ctx1;
wire MEMC73_write_mem_en_ctx1;
wire MEMC73_mem_en_ctx1;
wire [5:0] MEMC73_start_addr_ctx1;
wire [0:0] MEMC73_stride_ctx1;
wire [5:0] MEMC73_addr_out_ctx2;
wire MEMC73_write_en_ctx2;
wire MEMC73_write_mem_en_ctx2;
wire MEMC73_mem_en_ctx2;
wire [5:0] MEMC73_start_addr_ctx2;
wire [0:0] MEMC73_stride_ctx2;
wire [31:0] MEMC73_data_in_ctx1;
wire [31:0] MEMC73_data_in_ctx2;
wire [31:0] MEMC73_data_out_ctx1;
wire [31:0] MEMC73_data_out_ctx2;
wire [63:0] MEMC73_burst_count_ctx1;
wire [63:0] MEMC73_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC73(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC73_data_from_Core),
.data_to_Core(MEMC73_data_to_Core),
.valid_ctx1(MEMC73_valid_ctx1),
.addr_out_ctx1(MEMC73_addr_out_ctx1),
.write_en_ctx1(MEMC73_write_en_ctx1),
.start_addr_ctx1(MEMC73_start_addr_ctx1),
.stride_ctx1(MEMC73_stride_ctx1),
.burst_count_ctx1(MEMC73_burst_count_ctx1),
.valid_ctx2(MEMC73_valid_ctx2),
.addr_out_ctx2(MEMC73_addr_out_ctx2),
.write_en_ctx2(MEMC73_write_en_ctx2),
.start_addr_ctx2(MEMC73_start_addr_ctx2),
.stride_ctx2(MEMC73_stride_ctx2),
.burst_count_ctx2(MEMC73_burst_count_ctx2),
.data_in_ctx1(MEMC73_data_in_ctx1),
.data_in_ctx2(MEMC73_data_in_ctx2),
.data_out_ctx1(MEMC73_data_out_ctx1),
.data_out_ctx2(MEMC73_data_out_ctx2),
.write_mem_en_ctx1(MEMC73_write_mem_en_ctx1),
.mem_en_ctx1(MEMC73_mem_en_ctx1),.write_mem_en_ctx2(MEMC73_write_mem_en_ctx2),
.mem_en_ctx2(MEMC73_mem_en_ctx2));

defparam MEMC73.DATA_WIDTH = 32;
defparam MEMC73.ADDR_WIDTH = 6;
defparam MEMC73.STRIDE_WIDTH = 1;
wire MEMC74_valid_ctx1;
wire MEMC74_valid_ctx2;
wire [31:0] MEMC74_data_from_Core;
wire [31:0] MEMC74_data_to_Core;
wire [5:0] MEMC74_addr_out_ctx1;
wire MEMC74_write_en_ctx1;
wire MEMC74_write_mem_en_ctx1;
wire MEMC74_mem_en_ctx1;
wire [5:0] MEMC74_start_addr_ctx1;
wire [0:0] MEMC74_stride_ctx1;
wire [5:0] MEMC74_addr_out_ctx2;
wire MEMC74_write_en_ctx2;
wire MEMC74_write_mem_en_ctx2;
wire MEMC74_mem_en_ctx2;
wire [5:0] MEMC74_start_addr_ctx2;
wire [0:0] MEMC74_stride_ctx2;
wire [31:0] MEMC74_data_in_ctx1;
wire [31:0] MEMC74_data_in_ctx2;
wire [31:0] MEMC74_data_out_ctx1;
wire [31:0] MEMC74_data_out_ctx2;
wire [63:0] MEMC74_burst_count_ctx1;
wire [63:0] MEMC74_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC74(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC74_data_from_Core),
.data_to_Core(MEMC74_data_to_Core),
.valid_ctx1(MEMC74_valid_ctx1),
.addr_out_ctx1(MEMC74_addr_out_ctx1),
.write_en_ctx1(MEMC74_write_en_ctx1),
.start_addr_ctx1(MEMC74_start_addr_ctx1),
.stride_ctx1(MEMC74_stride_ctx1),
.burst_count_ctx1(MEMC74_burst_count_ctx1),
.valid_ctx2(MEMC74_valid_ctx2),
.addr_out_ctx2(MEMC74_addr_out_ctx2),
.write_en_ctx2(MEMC74_write_en_ctx2),
.start_addr_ctx2(MEMC74_start_addr_ctx2),
.stride_ctx2(MEMC74_stride_ctx2),
.burst_count_ctx2(MEMC74_burst_count_ctx2),
.data_in_ctx1(MEMC74_data_in_ctx1),
.data_in_ctx2(MEMC74_data_in_ctx2),
.data_out_ctx1(MEMC74_data_out_ctx1),
.data_out_ctx2(MEMC74_data_out_ctx2),
.write_mem_en_ctx1(MEMC74_write_mem_en_ctx1),
.mem_en_ctx1(MEMC74_mem_en_ctx1),.write_mem_en_ctx2(MEMC74_write_mem_en_ctx2),
.mem_en_ctx2(MEMC74_mem_en_ctx2));

defparam MEMC74.DATA_WIDTH = 32;
defparam MEMC74.ADDR_WIDTH = 6;
defparam MEMC74.STRIDE_WIDTH = 1;
wire MEMC75_valid_ctx1;
wire MEMC75_valid_ctx2;
wire [31:0] MEMC75_data_from_Core;
wire [31:0] MEMC75_data_to_Core;
wire [5:0] MEMC75_addr_out_ctx1;
wire MEMC75_write_en_ctx1;
wire MEMC75_write_mem_en_ctx1;
wire MEMC75_mem_en_ctx1;
wire [5:0] MEMC75_start_addr_ctx1;
wire [0:0] MEMC75_stride_ctx1;
wire [5:0] MEMC75_addr_out_ctx2;
wire MEMC75_write_en_ctx2;
wire MEMC75_write_mem_en_ctx2;
wire MEMC75_mem_en_ctx2;
wire [5:0] MEMC75_start_addr_ctx2;
wire [0:0] MEMC75_stride_ctx2;
wire [31:0] MEMC75_data_in_ctx1;
wire [31:0] MEMC75_data_in_ctx2;
wire [31:0] MEMC75_data_out_ctx1;
wire [31:0] MEMC75_data_out_ctx2;
wire [63:0] MEMC75_burst_count_ctx1;
wire [63:0] MEMC75_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC75(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC75_data_from_Core),
.data_to_Core(MEMC75_data_to_Core),
.valid_ctx1(MEMC75_valid_ctx1),
.addr_out_ctx1(MEMC75_addr_out_ctx1),
.write_en_ctx1(MEMC75_write_en_ctx1),
.start_addr_ctx1(MEMC75_start_addr_ctx1),
.stride_ctx1(MEMC75_stride_ctx1),
.burst_count_ctx1(MEMC75_burst_count_ctx1),
.valid_ctx2(MEMC75_valid_ctx2),
.addr_out_ctx2(MEMC75_addr_out_ctx2),
.write_en_ctx2(MEMC75_write_en_ctx2),
.start_addr_ctx2(MEMC75_start_addr_ctx2),
.stride_ctx2(MEMC75_stride_ctx2),
.burst_count_ctx2(MEMC75_burst_count_ctx2),
.data_in_ctx1(MEMC75_data_in_ctx1),
.data_in_ctx2(MEMC75_data_in_ctx2),
.data_out_ctx1(MEMC75_data_out_ctx1),
.data_out_ctx2(MEMC75_data_out_ctx2),
.write_mem_en_ctx1(MEMC75_write_mem_en_ctx1),
.mem_en_ctx1(MEMC75_mem_en_ctx1),.write_mem_en_ctx2(MEMC75_write_mem_en_ctx2),
.mem_en_ctx2(MEMC75_mem_en_ctx2));

defparam MEMC75.DATA_WIDTH = 32;
defparam MEMC75.ADDR_WIDTH = 6;
defparam MEMC75.STRIDE_WIDTH = 1;
wire MEMC76_valid_ctx1;
wire MEMC76_valid_ctx2;
wire [31:0] MEMC76_data_from_Core;
wire [31:0] MEMC76_data_to_Core;
wire [5:0] MEMC76_addr_out_ctx1;
wire MEMC76_write_en_ctx1;
wire MEMC76_write_mem_en_ctx1;
wire MEMC76_mem_en_ctx1;
wire [5:0] MEMC76_start_addr_ctx1;
wire [0:0] MEMC76_stride_ctx1;
wire [5:0] MEMC76_addr_out_ctx2;
wire MEMC76_write_en_ctx2;
wire MEMC76_write_mem_en_ctx2;
wire MEMC76_mem_en_ctx2;
wire [5:0] MEMC76_start_addr_ctx2;
wire [0:0] MEMC76_stride_ctx2;
wire [31:0] MEMC76_data_in_ctx1;
wire [31:0] MEMC76_data_in_ctx2;
wire [31:0] MEMC76_data_out_ctx1;
wire [31:0] MEMC76_data_out_ctx2;
wire [63:0] MEMC76_burst_count_ctx1;
wire [63:0] MEMC76_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC76(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC76_data_from_Core),
.data_to_Core(MEMC76_data_to_Core),
.valid_ctx1(MEMC76_valid_ctx1),
.addr_out_ctx1(MEMC76_addr_out_ctx1),
.write_en_ctx1(MEMC76_write_en_ctx1),
.start_addr_ctx1(MEMC76_start_addr_ctx1),
.stride_ctx1(MEMC76_stride_ctx1),
.burst_count_ctx1(MEMC76_burst_count_ctx1),
.valid_ctx2(MEMC76_valid_ctx2),
.addr_out_ctx2(MEMC76_addr_out_ctx2),
.write_en_ctx2(MEMC76_write_en_ctx2),
.start_addr_ctx2(MEMC76_start_addr_ctx2),
.stride_ctx2(MEMC76_stride_ctx2),
.burst_count_ctx2(MEMC76_burst_count_ctx2),
.data_in_ctx1(MEMC76_data_in_ctx1),
.data_in_ctx2(MEMC76_data_in_ctx2),
.data_out_ctx1(MEMC76_data_out_ctx1),
.data_out_ctx2(MEMC76_data_out_ctx2),
.write_mem_en_ctx1(MEMC76_write_mem_en_ctx1),
.mem_en_ctx1(MEMC76_mem_en_ctx1),.write_mem_en_ctx2(MEMC76_write_mem_en_ctx2),
.mem_en_ctx2(MEMC76_mem_en_ctx2));

defparam MEMC76.DATA_WIDTH = 32;
defparam MEMC76.ADDR_WIDTH = 6;
defparam MEMC76.STRIDE_WIDTH = 1;
wire MEMC77_valid_ctx1;
wire MEMC77_valid_ctx2;
wire [31:0] MEMC77_data_from_Core;
wire [31:0] MEMC77_data_to_Core;
wire [5:0] MEMC77_addr_out_ctx1;
wire MEMC77_write_en_ctx1;
wire MEMC77_write_mem_en_ctx1;
wire MEMC77_mem_en_ctx1;
wire [5:0] MEMC77_start_addr_ctx1;
wire [0:0] MEMC77_stride_ctx1;
wire [5:0] MEMC77_addr_out_ctx2;
wire MEMC77_write_en_ctx2;
wire MEMC77_write_mem_en_ctx2;
wire MEMC77_mem_en_ctx2;
wire [5:0] MEMC77_start_addr_ctx2;
wire [0:0] MEMC77_stride_ctx2;
wire [31:0] MEMC77_data_in_ctx1;
wire [31:0] MEMC77_data_in_ctx2;
wire [31:0] MEMC77_data_out_ctx1;
wire [31:0] MEMC77_data_out_ctx2;
wire [63:0] MEMC77_burst_count_ctx1;
wire [63:0] MEMC77_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC77(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC77_data_from_Core),
.data_to_Core(MEMC77_data_to_Core),
.valid_ctx1(MEMC77_valid_ctx1),
.addr_out_ctx1(MEMC77_addr_out_ctx1),
.write_en_ctx1(MEMC77_write_en_ctx1),
.start_addr_ctx1(MEMC77_start_addr_ctx1),
.stride_ctx1(MEMC77_stride_ctx1),
.burst_count_ctx1(MEMC77_burst_count_ctx1),
.valid_ctx2(MEMC77_valid_ctx2),
.addr_out_ctx2(MEMC77_addr_out_ctx2),
.write_en_ctx2(MEMC77_write_en_ctx2),
.start_addr_ctx2(MEMC77_start_addr_ctx2),
.stride_ctx2(MEMC77_stride_ctx2),
.burst_count_ctx2(MEMC77_burst_count_ctx2),
.data_in_ctx1(MEMC77_data_in_ctx1),
.data_in_ctx2(MEMC77_data_in_ctx2),
.data_out_ctx1(MEMC77_data_out_ctx1),
.data_out_ctx2(MEMC77_data_out_ctx2),
.write_mem_en_ctx1(MEMC77_write_mem_en_ctx1),
.mem_en_ctx1(MEMC77_mem_en_ctx1),.write_mem_en_ctx2(MEMC77_write_mem_en_ctx2),
.mem_en_ctx2(MEMC77_mem_en_ctx2));

defparam MEMC77.DATA_WIDTH = 32;
defparam MEMC77.ADDR_WIDTH = 6;
defparam MEMC77.STRIDE_WIDTH = 1;
wire MEMC78_valid_ctx1;
wire MEMC78_valid_ctx2;
wire [31:0] MEMC78_data_from_Core;
wire [31:0] MEMC78_data_to_Core;
wire [5:0] MEMC78_addr_out_ctx1;
wire MEMC78_write_en_ctx1;
wire MEMC78_write_mem_en_ctx1;
wire MEMC78_mem_en_ctx1;
wire [5:0] MEMC78_start_addr_ctx1;
wire [0:0] MEMC78_stride_ctx1;
wire [5:0] MEMC78_addr_out_ctx2;
wire MEMC78_write_en_ctx2;
wire MEMC78_write_mem_en_ctx2;
wire MEMC78_mem_en_ctx2;
wire [5:0] MEMC78_start_addr_ctx2;
wire [0:0] MEMC78_stride_ctx2;
wire [31:0] MEMC78_data_in_ctx1;
wire [31:0] MEMC78_data_in_ctx2;
wire [31:0] MEMC78_data_out_ctx1;
wire [31:0] MEMC78_data_out_ctx2;
wire [63:0] MEMC78_burst_count_ctx1;
wire [63:0] MEMC78_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC78(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC78_data_from_Core),
.data_to_Core(MEMC78_data_to_Core),
.valid_ctx1(MEMC78_valid_ctx1),
.addr_out_ctx1(MEMC78_addr_out_ctx1),
.write_en_ctx1(MEMC78_write_en_ctx1),
.start_addr_ctx1(MEMC78_start_addr_ctx1),
.stride_ctx1(MEMC78_stride_ctx1),
.burst_count_ctx1(MEMC78_burst_count_ctx1),
.valid_ctx2(MEMC78_valid_ctx2),
.addr_out_ctx2(MEMC78_addr_out_ctx2),
.write_en_ctx2(MEMC78_write_en_ctx2),
.start_addr_ctx2(MEMC78_start_addr_ctx2),
.stride_ctx2(MEMC78_stride_ctx2),
.burst_count_ctx2(MEMC78_burst_count_ctx2),
.data_in_ctx1(MEMC78_data_in_ctx1),
.data_in_ctx2(MEMC78_data_in_ctx2),
.data_out_ctx1(MEMC78_data_out_ctx1),
.data_out_ctx2(MEMC78_data_out_ctx2),
.write_mem_en_ctx1(MEMC78_write_mem_en_ctx1),
.mem_en_ctx1(MEMC78_mem_en_ctx1),.write_mem_en_ctx2(MEMC78_write_mem_en_ctx2),
.mem_en_ctx2(MEMC78_mem_en_ctx2));

defparam MEMC78.DATA_WIDTH = 32;
defparam MEMC78.ADDR_WIDTH = 6;
defparam MEMC78.STRIDE_WIDTH = 1;
wire MEMC79_valid_ctx1;
wire MEMC79_valid_ctx2;
wire [31:0] MEMC79_data_from_Core;
wire [31:0] MEMC79_data_to_Core;
wire [5:0] MEMC79_addr_out_ctx1;
wire MEMC79_write_en_ctx1;
wire MEMC79_write_mem_en_ctx1;
wire MEMC79_mem_en_ctx1;
wire [5:0] MEMC79_start_addr_ctx1;
wire [0:0] MEMC79_stride_ctx1;
wire [5:0] MEMC79_addr_out_ctx2;
wire MEMC79_write_en_ctx2;
wire MEMC79_write_mem_en_ctx2;
wire MEMC79_mem_en_ctx2;
wire [5:0] MEMC79_start_addr_ctx2;
wire [0:0] MEMC79_stride_ctx2;
wire [31:0] MEMC79_data_in_ctx1;
wire [31:0] MEMC79_data_in_ctx2;
wire [31:0] MEMC79_data_out_ctx1;
wire [31:0] MEMC79_data_out_ctx2;
wire [63:0] MEMC79_burst_count_ctx1;
wire [63:0] MEMC79_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC79(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC79_data_from_Core),
.data_to_Core(MEMC79_data_to_Core),
.valid_ctx1(MEMC79_valid_ctx1),
.addr_out_ctx1(MEMC79_addr_out_ctx1),
.write_en_ctx1(MEMC79_write_en_ctx1),
.start_addr_ctx1(MEMC79_start_addr_ctx1),
.stride_ctx1(MEMC79_stride_ctx1),
.burst_count_ctx1(MEMC79_burst_count_ctx1),
.valid_ctx2(MEMC79_valid_ctx2),
.addr_out_ctx2(MEMC79_addr_out_ctx2),
.write_en_ctx2(MEMC79_write_en_ctx2),
.start_addr_ctx2(MEMC79_start_addr_ctx2),
.stride_ctx2(MEMC79_stride_ctx2),
.burst_count_ctx2(MEMC79_burst_count_ctx2),
.data_in_ctx1(MEMC79_data_in_ctx1),
.data_in_ctx2(MEMC79_data_in_ctx2),
.data_out_ctx1(MEMC79_data_out_ctx1),
.data_out_ctx2(MEMC79_data_out_ctx2),
.write_mem_en_ctx1(MEMC79_write_mem_en_ctx1),
.mem_en_ctx1(MEMC79_mem_en_ctx1),.write_mem_en_ctx2(MEMC79_write_mem_en_ctx2),
.mem_en_ctx2(MEMC79_mem_en_ctx2));

defparam MEMC79.DATA_WIDTH = 32;
defparam MEMC79.ADDR_WIDTH = 6;
defparam MEMC79.STRIDE_WIDTH = 1;
wire MEMC80_valid_ctx1;
wire MEMC80_valid_ctx2;
wire [31:0] MEMC80_data_from_Core;
wire [31:0] MEMC80_data_to_Core;
wire [5:0] MEMC80_addr_out_ctx1;
wire MEMC80_write_en_ctx1;
wire MEMC80_write_mem_en_ctx1;
wire MEMC80_mem_en_ctx1;
wire [5:0] MEMC80_start_addr_ctx1;
wire [0:0] MEMC80_stride_ctx1;
wire [5:0] MEMC80_addr_out_ctx2;
wire MEMC80_write_en_ctx2;
wire MEMC80_write_mem_en_ctx2;
wire MEMC80_mem_en_ctx2;
wire [5:0] MEMC80_start_addr_ctx2;
wire [0:0] MEMC80_stride_ctx2;
wire [31:0] MEMC80_data_in_ctx1;
wire [31:0] MEMC80_data_in_ctx2;
wire [31:0] MEMC80_data_out_ctx1;
wire [31:0] MEMC80_data_out_ctx2;
wire [63:0] MEMC80_burst_count_ctx1;
wire [63:0] MEMC80_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC80(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC80_data_from_Core),
.data_to_Core(MEMC80_data_to_Core),
.valid_ctx1(MEMC80_valid_ctx1),
.addr_out_ctx1(MEMC80_addr_out_ctx1),
.write_en_ctx1(MEMC80_write_en_ctx1),
.start_addr_ctx1(MEMC80_start_addr_ctx1),
.stride_ctx1(MEMC80_stride_ctx1),
.burst_count_ctx1(MEMC80_burst_count_ctx1),
.valid_ctx2(MEMC80_valid_ctx2),
.addr_out_ctx2(MEMC80_addr_out_ctx2),
.write_en_ctx2(MEMC80_write_en_ctx2),
.start_addr_ctx2(MEMC80_start_addr_ctx2),
.stride_ctx2(MEMC80_stride_ctx2),
.burst_count_ctx2(MEMC80_burst_count_ctx2),
.data_in_ctx1(MEMC80_data_in_ctx1),
.data_in_ctx2(MEMC80_data_in_ctx2),
.data_out_ctx1(MEMC80_data_out_ctx1),
.data_out_ctx2(MEMC80_data_out_ctx2),
.write_mem_en_ctx1(MEMC80_write_mem_en_ctx1),
.mem_en_ctx1(MEMC80_mem_en_ctx1),.write_mem_en_ctx2(MEMC80_write_mem_en_ctx2),
.mem_en_ctx2(MEMC80_mem_en_ctx2));

defparam MEMC80.DATA_WIDTH = 32;
defparam MEMC80.ADDR_WIDTH = 6;
defparam MEMC80.STRIDE_WIDTH = 1;
wire MEMC81_valid_ctx1;
wire MEMC81_valid_ctx2;
wire [31:0] MEMC81_data_from_Core;
wire [31:0] MEMC81_data_to_Core;
wire [5:0] MEMC81_addr_out_ctx1;
wire MEMC81_write_en_ctx1;
wire MEMC81_write_mem_en_ctx1;
wire MEMC81_mem_en_ctx1;
wire [5:0] MEMC81_start_addr_ctx1;
wire [0:0] MEMC81_stride_ctx1;
wire [5:0] MEMC81_addr_out_ctx2;
wire MEMC81_write_en_ctx2;
wire MEMC81_write_mem_en_ctx2;
wire MEMC81_mem_en_ctx2;
wire [5:0] MEMC81_start_addr_ctx2;
wire [0:0] MEMC81_stride_ctx2;
wire [31:0] MEMC81_data_in_ctx1;
wire [31:0] MEMC81_data_in_ctx2;
wire [31:0] MEMC81_data_out_ctx1;
wire [31:0] MEMC81_data_out_ctx2;
wire [63:0] MEMC81_burst_count_ctx1;
wire [63:0] MEMC81_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC81(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC81_data_from_Core),
.data_to_Core(MEMC81_data_to_Core),
.valid_ctx1(MEMC81_valid_ctx1),
.addr_out_ctx1(MEMC81_addr_out_ctx1),
.write_en_ctx1(MEMC81_write_en_ctx1),
.start_addr_ctx1(MEMC81_start_addr_ctx1),
.stride_ctx1(MEMC81_stride_ctx1),
.burst_count_ctx1(MEMC81_burst_count_ctx1),
.valid_ctx2(MEMC81_valid_ctx2),
.addr_out_ctx2(MEMC81_addr_out_ctx2),
.write_en_ctx2(MEMC81_write_en_ctx2),
.start_addr_ctx2(MEMC81_start_addr_ctx2),
.stride_ctx2(MEMC81_stride_ctx2),
.burst_count_ctx2(MEMC81_burst_count_ctx2),
.data_in_ctx1(MEMC81_data_in_ctx1),
.data_in_ctx2(MEMC81_data_in_ctx2),
.data_out_ctx1(MEMC81_data_out_ctx1),
.data_out_ctx2(MEMC81_data_out_ctx2),
.write_mem_en_ctx1(MEMC81_write_mem_en_ctx1),
.mem_en_ctx1(MEMC81_mem_en_ctx1),.write_mem_en_ctx2(MEMC81_write_mem_en_ctx2),
.mem_en_ctx2(MEMC81_mem_en_ctx2));

defparam MEMC81.DATA_WIDTH = 32;
defparam MEMC81.ADDR_WIDTH = 6;
defparam MEMC81.STRIDE_WIDTH = 1;
wire MEMC82_valid_ctx1;
wire MEMC82_valid_ctx2;
wire [31:0] MEMC82_data_from_Core;
wire [31:0] MEMC82_data_to_Core;
wire [5:0] MEMC82_addr_out_ctx1;
wire MEMC82_write_en_ctx1;
wire MEMC82_write_mem_en_ctx1;
wire MEMC82_mem_en_ctx1;
wire [5:0] MEMC82_start_addr_ctx1;
wire [0:0] MEMC82_stride_ctx1;
wire [5:0] MEMC82_addr_out_ctx2;
wire MEMC82_write_en_ctx2;
wire MEMC82_write_mem_en_ctx2;
wire MEMC82_mem_en_ctx2;
wire [5:0] MEMC82_start_addr_ctx2;
wire [0:0] MEMC82_stride_ctx2;
wire [31:0] MEMC82_data_in_ctx1;
wire [31:0] MEMC82_data_in_ctx2;
wire [31:0] MEMC82_data_out_ctx1;
wire [31:0] MEMC82_data_out_ctx2;
wire [63:0] MEMC82_burst_count_ctx1;
wire [63:0] MEMC82_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC82(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC82_data_from_Core),
.data_to_Core(MEMC82_data_to_Core),
.valid_ctx1(MEMC82_valid_ctx1),
.addr_out_ctx1(MEMC82_addr_out_ctx1),
.write_en_ctx1(MEMC82_write_en_ctx1),
.start_addr_ctx1(MEMC82_start_addr_ctx1),
.stride_ctx1(MEMC82_stride_ctx1),
.burst_count_ctx1(MEMC82_burst_count_ctx1),
.valid_ctx2(MEMC82_valid_ctx2),
.addr_out_ctx2(MEMC82_addr_out_ctx2),
.write_en_ctx2(MEMC82_write_en_ctx2),
.start_addr_ctx2(MEMC82_start_addr_ctx2),
.stride_ctx2(MEMC82_stride_ctx2),
.burst_count_ctx2(MEMC82_burst_count_ctx2),
.data_in_ctx1(MEMC82_data_in_ctx1),
.data_in_ctx2(MEMC82_data_in_ctx2),
.data_out_ctx1(MEMC82_data_out_ctx1),
.data_out_ctx2(MEMC82_data_out_ctx2),
.write_mem_en_ctx1(MEMC82_write_mem_en_ctx1),
.mem_en_ctx1(MEMC82_mem_en_ctx1),.write_mem_en_ctx2(MEMC82_write_mem_en_ctx2),
.mem_en_ctx2(MEMC82_mem_en_ctx2));

defparam MEMC82.DATA_WIDTH = 32;
defparam MEMC82.ADDR_WIDTH = 6;
defparam MEMC82.STRIDE_WIDTH = 1;
wire MEMC83_valid_ctx1;
wire MEMC83_valid_ctx2;
wire [31:0] MEMC83_data_from_Core;
wire [31:0] MEMC83_data_to_Core;
wire [5:0] MEMC83_addr_out_ctx1;
wire MEMC83_write_en_ctx1;
wire MEMC83_write_mem_en_ctx1;
wire MEMC83_mem_en_ctx1;
wire [5:0] MEMC83_start_addr_ctx1;
wire [0:0] MEMC83_stride_ctx1;
wire [5:0] MEMC83_addr_out_ctx2;
wire MEMC83_write_en_ctx2;
wire MEMC83_write_mem_en_ctx2;
wire MEMC83_mem_en_ctx2;
wire [5:0] MEMC83_start_addr_ctx2;
wire [0:0] MEMC83_stride_ctx2;
wire [31:0] MEMC83_data_in_ctx1;
wire [31:0] MEMC83_data_in_ctx2;
wire [31:0] MEMC83_data_out_ctx1;
wire [31:0] MEMC83_data_out_ctx2;
wire [63:0] MEMC83_burst_count_ctx1;
wire [63:0] MEMC83_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC83(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC83_data_from_Core),
.data_to_Core(MEMC83_data_to_Core),
.valid_ctx1(MEMC83_valid_ctx1),
.addr_out_ctx1(MEMC83_addr_out_ctx1),
.write_en_ctx1(MEMC83_write_en_ctx1),
.start_addr_ctx1(MEMC83_start_addr_ctx1),
.stride_ctx1(MEMC83_stride_ctx1),
.burst_count_ctx1(MEMC83_burst_count_ctx1),
.valid_ctx2(MEMC83_valid_ctx2),
.addr_out_ctx2(MEMC83_addr_out_ctx2),
.write_en_ctx2(MEMC83_write_en_ctx2),
.start_addr_ctx2(MEMC83_start_addr_ctx2),
.stride_ctx2(MEMC83_stride_ctx2),
.burst_count_ctx2(MEMC83_burst_count_ctx2),
.data_in_ctx1(MEMC83_data_in_ctx1),
.data_in_ctx2(MEMC83_data_in_ctx2),
.data_out_ctx1(MEMC83_data_out_ctx1),
.data_out_ctx2(MEMC83_data_out_ctx2),
.write_mem_en_ctx1(MEMC83_write_mem_en_ctx1),
.mem_en_ctx1(MEMC83_mem_en_ctx1),.write_mem_en_ctx2(MEMC83_write_mem_en_ctx2),
.mem_en_ctx2(MEMC83_mem_en_ctx2));

defparam MEMC83.DATA_WIDTH = 32;
defparam MEMC83.ADDR_WIDTH = 6;
defparam MEMC83.STRIDE_WIDTH = 1;
wire MEMC84_valid_ctx1;
wire MEMC84_valid_ctx2;
wire [31:0] MEMC84_data_from_Core;
wire [31:0] MEMC84_data_to_Core;
wire [5:0] MEMC84_addr_out_ctx1;
wire MEMC84_write_en_ctx1;
wire MEMC84_write_mem_en_ctx1;
wire MEMC84_mem_en_ctx1;
wire [5:0] MEMC84_start_addr_ctx1;
wire [0:0] MEMC84_stride_ctx1;
wire [5:0] MEMC84_addr_out_ctx2;
wire MEMC84_write_en_ctx2;
wire MEMC84_write_mem_en_ctx2;
wire MEMC84_mem_en_ctx2;
wire [5:0] MEMC84_start_addr_ctx2;
wire [0:0] MEMC84_stride_ctx2;
wire [31:0] MEMC84_data_in_ctx1;
wire [31:0] MEMC84_data_in_ctx2;
wire [31:0] MEMC84_data_out_ctx1;
wire [31:0] MEMC84_data_out_ctx2;
wire [63:0] MEMC84_burst_count_ctx1;
wire [63:0] MEMC84_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC84(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC84_data_from_Core),
.data_to_Core(MEMC84_data_to_Core),
.valid_ctx1(MEMC84_valid_ctx1),
.addr_out_ctx1(MEMC84_addr_out_ctx1),
.write_en_ctx1(MEMC84_write_en_ctx1),
.start_addr_ctx1(MEMC84_start_addr_ctx1),
.stride_ctx1(MEMC84_stride_ctx1),
.burst_count_ctx1(MEMC84_burst_count_ctx1),
.valid_ctx2(MEMC84_valid_ctx2),
.addr_out_ctx2(MEMC84_addr_out_ctx2),
.write_en_ctx2(MEMC84_write_en_ctx2),
.start_addr_ctx2(MEMC84_start_addr_ctx2),
.stride_ctx2(MEMC84_stride_ctx2),
.burst_count_ctx2(MEMC84_burst_count_ctx2),
.data_in_ctx1(MEMC84_data_in_ctx1),
.data_in_ctx2(MEMC84_data_in_ctx2),
.data_out_ctx1(MEMC84_data_out_ctx1),
.data_out_ctx2(MEMC84_data_out_ctx2),
.write_mem_en_ctx1(MEMC84_write_mem_en_ctx1),
.mem_en_ctx1(MEMC84_mem_en_ctx1),.write_mem_en_ctx2(MEMC84_write_mem_en_ctx2),
.mem_en_ctx2(MEMC84_mem_en_ctx2));

defparam MEMC84.DATA_WIDTH = 32;
defparam MEMC84.ADDR_WIDTH = 6;
defparam MEMC84.STRIDE_WIDTH = 1;
wire MEMC85_valid_ctx1;
wire MEMC85_valid_ctx2;
wire [31:0] MEMC85_data_from_Core;
wire [31:0] MEMC85_data_to_Core;
wire [5:0] MEMC85_addr_out_ctx1;
wire MEMC85_write_en_ctx1;
wire MEMC85_write_mem_en_ctx1;
wire MEMC85_mem_en_ctx1;
wire [5:0] MEMC85_start_addr_ctx1;
wire [0:0] MEMC85_stride_ctx1;
wire [5:0] MEMC85_addr_out_ctx2;
wire MEMC85_write_en_ctx2;
wire MEMC85_write_mem_en_ctx2;
wire MEMC85_mem_en_ctx2;
wire [5:0] MEMC85_start_addr_ctx2;
wire [0:0] MEMC85_stride_ctx2;
wire [31:0] MEMC85_data_in_ctx1;
wire [31:0] MEMC85_data_in_ctx2;
wire [31:0] MEMC85_data_out_ctx1;
wire [31:0] MEMC85_data_out_ctx2;
wire [63:0] MEMC85_burst_count_ctx1;
wire [63:0] MEMC85_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC85(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC85_data_from_Core),
.data_to_Core(MEMC85_data_to_Core),
.valid_ctx1(MEMC85_valid_ctx1),
.addr_out_ctx1(MEMC85_addr_out_ctx1),
.write_en_ctx1(MEMC85_write_en_ctx1),
.start_addr_ctx1(MEMC85_start_addr_ctx1),
.stride_ctx1(MEMC85_stride_ctx1),
.burst_count_ctx1(MEMC85_burst_count_ctx1),
.valid_ctx2(MEMC85_valid_ctx2),
.addr_out_ctx2(MEMC85_addr_out_ctx2),
.write_en_ctx2(MEMC85_write_en_ctx2),
.start_addr_ctx2(MEMC85_start_addr_ctx2),
.stride_ctx2(MEMC85_stride_ctx2),
.burst_count_ctx2(MEMC85_burst_count_ctx2),
.data_in_ctx1(MEMC85_data_in_ctx1),
.data_in_ctx2(MEMC85_data_in_ctx2),
.data_out_ctx1(MEMC85_data_out_ctx1),
.data_out_ctx2(MEMC85_data_out_ctx2),
.write_mem_en_ctx1(MEMC85_write_mem_en_ctx1),
.mem_en_ctx1(MEMC85_mem_en_ctx1),.write_mem_en_ctx2(MEMC85_write_mem_en_ctx2),
.mem_en_ctx2(MEMC85_mem_en_ctx2));

defparam MEMC85.DATA_WIDTH = 32;
defparam MEMC85.ADDR_WIDTH = 6;
defparam MEMC85.STRIDE_WIDTH = 1;
wire MEMC86_valid_ctx1;
wire MEMC86_valid_ctx2;
wire [31:0] MEMC86_data_from_Core;
wire [31:0] MEMC86_data_to_Core;
wire [5:0] MEMC86_addr_out_ctx1;
wire MEMC86_write_en_ctx1;
wire MEMC86_write_mem_en_ctx1;
wire MEMC86_mem_en_ctx1;
wire [5:0] MEMC86_start_addr_ctx1;
wire [0:0] MEMC86_stride_ctx1;
wire [5:0] MEMC86_addr_out_ctx2;
wire MEMC86_write_en_ctx2;
wire MEMC86_write_mem_en_ctx2;
wire MEMC86_mem_en_ctx2;
wire [5:0] MEMC86_start_addr_ctx2;
wire [0:0] MEMC86_stride_ctx2;
wire [31:0] MEMC86_data_in_ctx1;
wire [31:0] MEMC86_data_in_ctx2;
wire [31:0] MEMC86_data_out_ctx1;
wire [31:0] MEMC86_data_out_ctx2;
wire [63:0] MEMC86_burst_count_ctx1;
wire [63:0] MEMC86_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC86(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC86_data_from_Core),
.data_to_Core(MEMC86_data_to_Core),
.valid_ctx1(MEMC86_valid_ctx1),
.addr_out_ctx1(MEMC86_addr_out_ctx1),
.write_en_ctx1(MEMC86_write_en_ctx1),
.start_addr_ctx1(MEMC86_start_addr_ctx1),
.stride_ctx1(MEMC86_stride_ctx1),
.burst_count_ctx1(MEMC86_burst_count_ctx1),
.valid_ctx2(MEMC86_valid_ctx2),
.addr_out_ctx2(MEMC86_addr_out_ctx2),
.write_en_ctx2(MEMC86_write_en_ctx2),
.start_addr_ctx2(MEMC86_start_addr_ctx2),
.stride_ctx2(MEMC86_stride_ctx2),
.burst_count_ctx2(MEMC86_burst_count_ctx2),
.data_in_ctx1(MEMC86_data_in_ctx1),
.data_in_ctx2(MEMC86_data_in_ctx2),
.data_out_ctx1(MEMC86_data_out_ctx1),
.data_out_ctx2(MEMC86_data_out_ctx2),
.write_mem_en_ctx1(MEMC86_write_mem_en_ctx1),
.mem_en_ctx1(MEMC86_mem_en_ctx1),.write_mem_en_ctx2(MEMC86_write_mem_en_ctx2),
.mem_en_ctx2(MEMC86_mem_en_ctx2));

defparam MEMC86.DATA_WIDTH = 32;
defparam MEMC86.ADDR_WIDTH = 6;
defparam MEMC86.STRIDE_WIDTH = 1;
wire MEMC87_valid_ctx1;
wire MEMC87_valid_ctx2;
wire [31:0] MEMC87_data_from_Core;
wire [31:0] MEMC87_data_to_Core;
wire [5:0] MEMC87_addr_out_ctx1;
wire MEMC87_write_en_ctx1;
wire MEMC87_write_mem_en_ctx1;
wire MEMC87_mem_en_ctx1;
wire [5:0] MEMC87_start_addr_ctx1;
wire [0:0] MEMC87_stride_ctx1;
wire [5:0] MEMC87_addr_out_ctx2;
wire MEMC87_write_en_ctx2;
wire MEMC87_write_mem_en_ctx2;
wire MEMC87_mem_en_ctx2;
wire [5:0] MEMC87_start_addr_ctx2;
wire [0:0] MEMC87_stride_ctx2;
wire [31:0] MEMC87_data_in_ctx1;
wire [31:0] MEMC87_data_in_ctx2;
wire [31:0] MEMC87_data_out_ctx1;
wire [31:0] MEMC87_data_out_ctx2;
wire [63:0] MEMC87_burst_count_ctx1;
wire [63:0] MEMC87_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC87(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC87_data_from_Core),
.data_to_Core(MEMC87_data_to_Core),
.valid_ctx1(MEMC87_valid_ctx1),
.addr_out_ctx1(MEMC87_addr_out_ctx1),
.write_en_ctx1(MEMC87_write_en_ctx1),
.start_addr_ctx1(MEMC87_start_addr_ctx1),
.stride_ctx1(MEMC87_stride_ctx1),
.burst_count_ctx1(MEMC87_burst_count_ctx1),
.valid_ctx2(MEMC87_valid_ctx2),
.addr_out_ctx2(MEMC87_addr_out_ctx2),
.write_en_ctx2(MEMC87_write_en_ctx2),
.start_addr_ctx2(MEMC87_start_addr_ctx2),
.stride_ctx2(MEMC87_stride_ctx2),
.burst_count_ctx2(MEMC87_burst_count_ctx2),
.data_in_ctx1(MEMC87_data_in_ctx1),
.data_in_ctx2(MEMC87_data_in_ctx2),
.data_out_ctx1(MEMC87_data_out_ctx1),
.data_out_ctx2(MEMC87_data_out_ctx2),
.write_mem_en_ctx1(MEMC87_write_mem_en_ctx1),
.mem_en_ctx1(MEMC87_mem_en_ctx1),.write_mem_en_ctx2(MEMC87_write_mem_en_ctx2),
.mem_en_ctx2(MEMC87_mem_en_ctx2));

defparam MEMC87.DATA_WIDTH = 32;
defparam MEMC87.ADDR_WIDTH = 6;
defparam MEMC87.STRIDE_WIDTH = 1;
wire MEMC88_valid_ctx1;
wire MEMC88_valid_ctx2;
wire [31:0] MEMC88_data_from_Core;
wire [31:0] MEMC88_data_to_Core;
wire [5:0] MEMC88_addr_out_ctx1;
wire MEMC88_write_en_ctx1;
wire MEMC88_write_mem_en_ctx1;
wire MEMC88_mem_en_ctx1;
wire [5:0] MEMC88_start_addr_ctx1;
wire [0:0] MEMC88_stride_ctx1;
wire [5:0] MEMC88_addr_out_ctx2;
wire MEMC88_write_en_ctx2;
wire MEMC88_write_mem_en_ctx2;
wire MEMC88_mem_en_ctx2;
wire [5:0] MEMC88_start_addr_ctx2;
wire [0:0] MEMC88_stride_ctx2;
wire [31:0] MEMC88_data_in_ctx1;
wire [31:0] MEMC88_data_in_ctx2;
wire [31:0] MEMC88_data_out_ctx1;
wire [31:0] MEMC88_data_out_ctx2;
wire [63:0] MEMC88_burst_count_ctx1;
wire [63:0] MEMC88_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC88(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC88_data_from_Core),
.data_to_Core(MEMC88_data_to_Core),
.valid_ctx1(MEMC88_valid_ctx1),
.addr_out_ctx1(MEMC88_addr_out_ctx1),
.write_en_ctx1(MEMC88_write_en_ctx1),
.start_addr_ctx1(MEMC88_start_addr_ctx1),
.stride_ctx1(MEMC88_stride_ctx1),
.burst_count_ctx1(MEMC88_burst_count_ctx1),
.valid_ctx2(MEMC88_valid_ctx2),
.addr_out_ctx2(MEMC88_addr_out_ctx2),
.write_en_ctx2(MEMC88_write_en_ctx2),
.start_addr_ctx2(MEMC88_start_addr_ctx2),
.stride_ctx2(MEMC88_stride_ctx2),
.burst_count_ctx2(MEMC88_burst_count_ctx2),
.data_in_ctx1(MEMC88_data_in_ctx1),
.data_in_ctx2(MEMC88_data_in_ctx2),
.data_out_ctx1(MEMC88_data_out_ctx1),
.data_out_ctx2(MEMC88_data_out_ctx2),
.write_mem_en_ctx1(MEMC88_write_mem_en_ctx1),
.mem_en_ctx1(MEMC88_mem_en_ctx1),.write_mem_en_ctx2(MEMC88_write_mem_en_ctx2),
.mem_en_ctx2(MEMC88_mem_en_ctx2));

defparam MEMC88.DATA_WIDTH = 32;
defparam MEMC88.ADDR_WIDTH = 6;
defparam MEMC88.STRIDE_WIDTH = 1;
wire MEMC89_valid_ctx1;
wire MEMC89_valid_ctx2;
wire [31:0] MEMC89_data_from_Core;
wire [31:0] MEMC89_data_to_Core;
wire [5:0] MEMC89_addr_out_ctx1;
wire MEMC89_write_en_ctx1;
wire MEMC89_write_mem_en_ctx1;
wire MEMC89_mem_en_ctx1;
wire [5:0] MEMC89_start_addr_ctx1;
wire [0:0] MEMC89_stride_ctx1;
wire [5:0] MEMC89_addr_out_ctx2;
wire MEMC89_write_en_ctx2;
wire MEMC89_write_mem_en_ctx2;
wire MEMC89_mem_en_ctx2;
wire [5:0] MEMC89_start_addr_ctx2;
wire [0:0] MEMC89_stride_ctx2;
wire [31:0] MEMC89_data_in_ctx1;
wire [31:0] MEMC89_data_in_ctx2;
wire [31:0] MEMC89_data_out_ctx1;
wire [31:0] MEMC89_data_out_ctx2;
wire [63:0] MEMC89_burst_count_ctx1;
wire [63:0] MEMC89_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC89(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC89_data_from_Core),
.data_to_Core(MEMC89_data_to_Core),
.valid_ctx1(MEMC89_valid_ctx1),
.addr_out_ctx1(MEMC89_addr_out_ctx1),
.write_en_ctx1(MEMC89_write_en_ctx1),
.start_addr_ctx1(MEMC89_start_addr_ctx1),
.stride_ctx1(MEMC89_stride_ctx1),
.burst_count_ctx1(MEMC89_burst_count_ctx1),
.valid_ctx2(MEMC89_valid_ctx2),
.addr_out_ctx2(MEMC89_addr_out_ctx2),
.write_en_ctx2(MEMC89_write_en_ctx2),
.start_addr_ctx2(MEMC89_start_addr_ctx2),
.stride_ctx2(MEMC89_stride_ctx2),
.burst_count_ctx2(MEMC89_burst_count_ctx2),
.data_in_ctx1(MEMC89_data_in_ctx1),
.data_in_ctx2(MEMC89_data_in_ctx2),
.data_out_ctx1(MEMC89_data_out_ctx1),
.data_out_ctx2(MEMC89_data_out_ctx2),
.write_mem_en_ctx1(MEMC89_write_mem_en_ctx1),
.mem_en_ctx1(MEMC89_mem_en_ctx1),.write_mem_en_ctx2(MEMC89_write_mem_en_ctx2),
.mem_en_ctx2(MEMC89_mem_en_ctx2));

defparam MEMC89.DATA_WIDTH = 32;
defparam MEMC89.ADDR_WIDTH = 6;
defparam MEMC89.STRIDE_WIDTH = 1;
wire MEMC90_valid_ctx1;
wire MEMC90_valid_ctx2;
wire [31:0] MEMC90_data_from_Core;
wire [31:0] MEMC90_data_to_Core;
wire [5:0] MEMC90_addr_out_ctx1;
wire MEMC90_write_en_ctx1;
wire MEMC90_write_mem_en_ctx1;
wire MEMC90_mem_en_ctx1;
wire [5:0] MEMC90_start_addr_ctx1;
wire [0:0] MEMC90_stride_ctx1;
wire [5:0] MEMC90_addr_out_ctx2;
wire MEMC90_write_en_ctx2;
wire MEMC90_write_mem_en_ctx2;
wire MEMC90_mem_en_ctx2;
wire [5:0] MEMC90_start_addr_ctx2;
wire [0:0] MEMC90_stride_ctx2;
wire [31:0] MEMC90_data_in_ctx1;
wire [31:0] MEMC90_data_in_ctx2;
wire [31:0] MEMC90_data_out_ctx1;
wire [31:0] MEMC90_data_out_ctx2;
wire [63:0] MEMC90_burst_count_ctx1;
wire [63:0] MEMC90_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC90(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC90_data_from_Core),
.data_to_Core(MEMC90_data_to_Core),
.valid_ctx1(MEMC90_valid_ctx1),
.addr_out_ctx1(MEMC90_addr_out_ctx1),
.write_en_ctx1(MEMC90_write_en_ctx1),
.start_addr_ctx1(MEMC90_start_addr_ctx1),
.stride_ctx1(MEMC90_stride_ctx1),
.burst_count_ctx1(MEMC90_burst_count_ctx1),
.valid_ctx2(MEMC90_valid_ctx2),
.addr_out_ctx2(MEMC90_addr_out_ctx2),
.write_en_ctx2(MEMC90_write_en_ctx2),
.start_addr_ctx2(MEMC90_start_addr_ctx2),
.stride_ctx2(MEMC90_stride_ctx2),
.burst_count_ctx2(MEMC90_burst_count_ctx2),
.data_in_ctx1(MEMC90_data_in_ctx1),
.data_in_ctx2(MEMC90_data_in_ctx2),
.data_out_ctx1(MEMC90_data_out_ctx1),
.data_out_ctx2(MEMC90_data_out_ctx2),
.write_mem_en_ctx1(MEMC90_write_mem_en_ctx1),
.mem_en_ctx1(MEMC90_mem_en_ctx1),.write_mem_en_ctx2(MEMC90_write_mem_en_ctx2),
.mem_en_ctx2(MEMC90_mem_en_ctx2));

defparam MEMC90.DATA_WIDTH = 32;
defparam MEMC90.ADDR_WIDTH = 6;
defparam MEMC90.STRIDE_WIDTH = 1;
wire MEMC91_valid_ctx1;
wire MEMC91_valid_ctx2;
wire [31:0] MEMC91_data_from_Core;
wire [31:0] MEMC91_data_to_Core;
wire [5:0] MEMC91_addr_out_ctx1;
wire MEMC91_write_en_ctx1;
wire MEMC91_write_mem_en_ctx1;
wire MEMC91_mem_en_ctx1;
wire [5:0] MEMC91_start_addr_ctx1;
wire [0:0] MEMC91_stride_ctx1;
wire [5:0] MEMC91_addr_out_ctx2;
wire MEMC91_write_en_ctx2;
wire MEMC91_write_mem_en_ctx2;
wire MEMC91_mem_en_ctx2;
wire [5:0] MEMC91_start_addr_ctx2;
wire [0:0] MEMC91_stride_ctx2;
wire [31:0] MEMC91_data_in_ctx1;
wire [31:0] MEMC91_data_in_ctx2;
wire [31:0] MEMC91_data_out_ctx1;
wire [31:0] MEMC91_data_out_ctx2;
wire [63:0] MEMC91_burst_count_ctx1;
wire [63:0] MEMC91_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC91(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC91_data_from_Core),
.data_to_Core(MEMC91_data_to_Core),
.valid_ctx1(MEMC91_valid_ctx1),
.addr_out_ctx1(MEMC91_addr_out_ctx1),
.write_en_ctx1(MEMC91_write_en_ctx1),
.start_addr_ctx1(MEMC91_start_addr_ctx1),
.stride_ctx1(MEMC91_stride_ctx1),
.burst_count_ctx1(MEMC91_burst_count_ctx1),
.valid_ctx2(MEMC91_valid_ctx2),
.addr_out_ctx2(MEMC91_addr_out_ctx2),
.write_en_ctx2(MEMC91_write_en_ctx2),
.start_addr_ctx2(MEMC91_start_addr_ctx2),
.stride_ctx2(MEMC91_stride_ctx2),
.burst_count_ctx2(MEMC91_burst_count_ctx2),
.data_in_ctx1(MEMC91_data_in_ctx1),
.data_in_ctx2(MEMC91_data_in_ctx2),
.data_out_ctx1(MEMC91_data_out_ctx1),
.data_out_ctx2(MEMC91_data_out_ctx2),
.write_mem_en_ctx1(MEMC91_write_mem_en_ctx1),
.mem_en_ctx1(MEMC91_mem_en_ctx1),.write_mem_en_ctx2(MEMC91_write_mem_en_ctx2),
.mem_en_ctx2(MEMC91_mem_en_ctx2));

defparam MEMC91.DATA_WIDTH = 32;
defparam MEMC91.ADDR_WIDTH = 6;
defparam MEMC91.STRIDE_WIDTH = 1;
wire MEMC92_valid_ctx1;
wire MEMC92_valid_ctx2;
wire [31:0] MEMC92_data_from_Core;
wire [31:0] MEMC92_data_to_Core;
wire [5:0] MEMC92_addr_out_ctx1;
wire MEMC92_write_en_ctx1;
wire MEMC92_write_mem_en_ctx1;
wire MEMC92_mem_en_ctx1;
wire [5:0] MEMC92_start_addr_ctx1;
wire [0:0] MEMC92_stride_ctx1;
wire [5:0] MEMC92_addr_out_ctx2;
wire MEMC92_write_en_ctx2;
wire MEMC92_write_mem_en_ctx2;
wire MEMC92_mem_en_ctx2;
wire [5:0] MEMC92_start_addr_ctx2;
wire [0:0] MEMC92_stride_ctx2;
wire [31:0] MEMC92_data_in_ctx1;
wire [31:0] MEMC92_data_in_ctx2;
wire [31:0] MEMC92_data_out_ctx1;
wire [31:0] MEMC92_data_out_ctx2;
wire [63:0] MEMC92_burst_count_ctx1;
wire [63:0] MEMC92_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC92(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC92_data_from_Core),
.data_to_Core(MEMC92_data_to_Core),
.valid_ctx1(MEMC92_valid_ctx1),
.addr_out_ctx1(MEMC92_addr_out_ctx1),
.write_en_ctx1(MEMC92_write_en_ctx1),
.start_addr_ctx1(MEMC92_start_addr_ctx1),
.stride_ctx1(MEMC92_stride_ctx1),
.burst_count_ctx1(MEMC92_burst_count_ctx1),
.valid_ctx2(MEMC92_valid_ctx2),
.addr_out_ctx2(MEMC92_addr_out_ctx2),
.write_en_ctx2(MEMC92_write_en_ctx2),
.start_addr_ctx2(MEMC92_start_addr_ctx2),
.stride_ctx2(MEMC92_stride_ctx2),
.burst_count_ctx2(MEMC92_burst_count_ctx2),
.data_in_ctx1(MEMC92_data_in_ctx1),
.data_in_ctx2(MEMC92_data_in_ctx2),
.data_out_ctx1(MEMC92_data_out_ctx1),
.data_out_ctx2(MEMC92_data_out_ctx2),
.write_mem_en_ctx1(MEMC92_write_mem_en_ctx1),
.mem_en_ctx1(MEMC92_mem_en_ctx1),.write_mem_en_ctx2(MEMC92_write_mem_en_ctx2),
.mem_en_ctx2(MEMC92_mem_en_ctx2));

defparam MEMC92.DATA_WIDTH = 32;
defparam MEMC92.ADDR_WIDTH = 6;
defparam MEMC92.STRIDE_WIDTH = 1;
wire MEMC93_valid_ctx1;
wire MEMC93_valid_ctx2;
wire [31:0] MEMC93_data_from_Core;
wire [31:0] MEMC93_data_to_Core;
wire [5:0] MEMC93_addr_out_ctx1;
wire MEMC93_write_en_ctx1;
wire MEMC93_write_mem_en_ctx1;
wire MEMC93_mem_en_ctx1;
wire [5:0] MEMC93_start_addr_ctx1;
wire [0:0] MEMC93_stride_ctx1;
wire [5:0] MEMC93_addr_out_ctx2;
wire MEMC93_write_en_ctx2;
wire MEMC93_write_mem_en_ctx2;
wire MEMC93_mem_en_ctx2;
wire [5:0] MEMC93_start_addr_ctx2;
wire [0:0] MEMC93_stride_ctx2;
wire [31:0] MEMC93_data_in_ctx1;
wire [31:0] MEMC93_data_in_ctx2;
wire [31:0] MEMC93_data_out_ctx1;
wire [31:0] MEMC93_data_out_ctx2;
wire [63:0] MEMC93_burst_count_ctx1;
wire [63:0] MEMC93_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC93(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC93_data_from_Core),
.data_to_Core(MEMC93_data_to_Core),
.valid_ctx1(MEMC93_valid_ctx1),
.addr_out_ctx1(MEMC93_addr_out_ctx1),
.write_en_ctx1(MEMC93_write_en_ctx1),
.start_addr_ctx1(MEMC93_start_addr_ctx1),
.stride_ctx1(MEMC93_stride_ctx1),
.burst_count_ctx1(MEMC93_burst_count_ctx1),
.valid_ctx2(MEMC93_valid_ctx2),
.addr_out_ctx2(MEMC93_addr_out_ctx2),
.write_en_ctx2(MEMC93_write_en_ctx2),
.start_addr_ctx2(MEMC93_start_addr_ctx2),
.stride_ctx2(MEMC93_stride_ctx2),
.burst_count_ctx2(MEMC93_burst_count_ctx2),
.data_in_ctx1(MEMC93_data_in_ctx1),
.data_in_ctx2(MEMC93_data_in_ctx2),
.data_out_ctx1(MEMC93_data_out_ctx1),
.data_out_ctx2(MEMC93_data_out_ctx2),
.write_mem_en_ctx1(MEMC93_write_mem_en_ctx1),
.mem_en_ctx1(MEMC93_mem_en_ctx1),.write_mem_en_ctx2(MEMC93_write_mem_en_ctx2),
.mem_en_ctx2(MEMC93_mem_en_ctx2));

defparam MEMC93.DATA_WIDTH = 32;
defparam MEMC93.ADDR_WIDTH = 6;
defparam MEMC93.STRIDE_WIDTH = 1;
wire MEMC94_valid_ctx1;
wire MEMC94_valid_ctx2;
wire [31:0] MEMC94_data_from_Core;
wire [31:0] MEMC94_data_to_Core;
wire [5:0] MEMC94_addr_out_ctx1;
wire MEMC94_write_en_ctx1;
wire MEMC94_write_mem_en_ctx1;
wire MEMC94_mem_en_ctx1;
wire [5:0] MEMC94_start_addr_ctx1;
wire [0:0] MEMC94_stride_ctx1;
wire [5:0] MEMC94_addr_out_ctx2;
wire MEMC94_write_en_ctx2;
wire MEMC94_write_mem_en_ctx2;
wire MEMC94_mem_en_ctx2;
wire [5:0] MEMC94_start_addr_ctx2;
wire [0:0] MEMC94_stride_ctx2;
wire [31:0] MEMC94_data_in_ctx1;
wire [31:0] MEMC94_data_in_ctx2;
wire [31:0] MEMC94_data_out_ctx1;
wire [31:0] MEMC94_data_out_ctx2;
wire [63:0] MEMC94_burst_count_ctx1;
wire [63:0] MEMC94_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC94(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC94_data_from_Core),
.data_to_Core(MEMC94_data_to_Core),
.valid_ctx1(MEMC94_valid_ctx1),
.addr_out_ctx1(MEMC94_addr_out_ctx1),
.write_en_ctx1(MEMC94_write_en_ctx1),
.start_addr_ctx1(MEMC94_start_addr_ctx1),
.stride_ctx1(MEMC94_stride_ctx1),
.burst_count_ctx1(MEMC94_burst_count_ctx1),
.valid_ctx2(MEMC94_valid_ctx2),
.addr_out_ctx2(MEMC94_addr_out_ctx2),
.write_en_ctx2(MEMC94_write_en_ctx2),
.start_addr_ctx2(MEMC94_start_addr_ctx2),
.stride_ctx2(MEMC94_stride_ctx2),
.burst_count_ctx2(MEMC94_burst_count_ctx2),
.data_in_ctx1(MEMC94_data_in_ctx1),
.data_in_ctx2(MEMC94_data_in_ctx2),
.data_out_ctx1(MEMC94_data_out_ctx1),
.data_out_ctx2(MEMC94_data_out_ctx2),
.write_mem_en_ctx1(MEMC94_write_mem_en_ctx1),
.mem_en_ctx1(MEMC94_mem_en_ctx1),.write_mem_en_ctx2(MEMC94_write_mem_en_ctx2),
.mem_en_ctx2(MEMC94_mem_en_ctx2));

defparam MEMC94.DATA_WIDTH = 32;
defparam MEMC94.ADDR_WIDTH = 6;
defparam MEMC94.STRIDE_WIDTH = 1;
wire MEMC95_valid_ctx1;
wire MEMC95_valid_ctx2;
wire [31:0] MEMC95_data_from_Core;
wire [31:0] MEMC95_data_to_Core;
wire [5:0] MEMC95_addr_out_ctx1;
wire MEMC95_write_en_ctx1;
wire MEMC95_write_mem_en_ctx1;
wire MEMC95_mem_en_ctx1;
wire [5:0] MEMC95_start_addr_ctx1;
wire [0:0] MEMC95_stride_ctx1;
wire [5:0] MEMC95_addr_out_ctx2;
wire MEMC95_write_en_ctx2;
wire MEMC95_write_mem_en_ctx2;
wire MEMC95_mem_en_ctx2;
wire [5:0] MEMC95_start_addr_ctx2;
wire [0:0] MEMC95_stride_ctx2;
wire [31:0] MEMC95_data_in_ctx1;
wire [31:0] MEMC95_data_in_ctx2;
wire [31:0] MEMC95_data_out_ctx1;
wire [31:0] MEMC95_data_out_ctx2;
wire [63:0] MEMC95_burst_count_ctx1;
wire [63:0] MEMC95_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC95(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC95_data_from_Core),
.data_to_Core(MEMC95_data_to_Core),
.valid_ctx1(MEMC95_valid_ctx1),
.addr_out_ctx1(MEMC95_addr_out_ctx1),
.write_en_ctx1(MEMC95_write_en_ctx1),
.start_addr_ctx1(MEMC95_start_addr_ctx1),
.stride_ctx1(MEMC95_stride_ctx1),
.burst_count_ctx1(MEMC95_burst_count_ctx1),
.valid_ctx2(MEMC95_valid_ctx2),
.addr_out_ctx2(MEMC95_addr_out_ctx2),
.write_en_ctx2(MEMC95_write_en_ctx2),
.start_addr_ctx2(MEMC95_start_addr_ctx2),
.stride_ctx2(MEMC95_stride_ctx2),
.burst_count_ctx2(MEMC95_burst_count_ctx2),
.data_in_ctx1(MEMC95_data_in_ctx1),
.data_in_ctx2(MEMC95_data_in_ctx2),
.data_out_ctx1(MEMC95_data_out_ctx1),
.data_out_ctx2(MEMC95_data_out_ctx2),
.write_mem_en_ctx1(MEMC95_write_mem_en_ctx1),
.mem_en_ctx1(MEMC95_mem_en_ctx1),.write_mem_en_ctx2(MEMC95_write_mem_en_ctx2),
.mem_en_ctx2(MEMC95_mem_en_ctx2));

defparam MEMC95.DATA_WIDTH = 32;
defparam MEMC95.ADDR_WIDTH = 6;
defparam MEMC95.STRIDE_WIDTH = 1;
wire MEMC96_valid_ctx1;
wire MEMC96_valid_ctx2;
wire [31:0] MEMC96_data_from_Core;
wire [31:0] MEMC96_data_to_Core;
wire [5:0] MEMC96_addr_out_ctx1;
wire MEMC96_write_en_ctx1;
wire MEMC96_write_mem_en_ctx1;
wire MEMC96_mem_en_ctx1;
wire [5:0] MEMC96_start_addr_ctx1;
wire [0:0] MEMC96_stride_ctx1;
wire [5:0] MEMC96_addr_out_ctx2;
wire MEMC96_write_en_ctx2;
wire MEMC96_write_mem_en_ctx2;
wire MEMC96_mem_en_ctx2;
wire [5:0] MEMC96_start_addr_ctx2;
wire [0:0] MEMC96_stride_ctx2;
wire [31:0] MEMC96_data_in_ctx1;
wire [31:0] MEMC96_data_in_ctx2;
wire [31:0] MEMC96_data_out_ctx1;
wire [31:0] MEMC96_data_out_ctx2;
wire [63:0] MEMC96_burst_count_ctx1;
wire [63:0] MEMC96_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC96(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC96_data_from_Core),
.data_to_Core(MEMC96_data_to_Core),
.valid_ctx1(MEMC96_valid_ctx1),
.addr_out_ctx1(MEMC96_addr_out_ctx1),
.write_en_ctx1(MEMC96_write_en_ctx1),
.start_addr_ctx1(MEMC96_start_addr_ctx1),
.stride_ctx1(MEMC96_stride_ctx1),
.burst_count_ctx1(MEMC96_burst_count_ctx1),
.valid_ctx2(MEMC96_valid_ctx2),
.addr_out_ctx2(MEMC96_addr_out_ctx2),
.write_en_ctx2(MEMC96_write_en_ctx2),
.start_addr_ctx2(MEMC96_start_addr_ctx2),
.stride_ctx2(MEMC96_stride_ctx2),
.burst_count_ctx2(MEMC96_burst_count_ctx2),
.data_in_ctx1(MEMC96_data_in_ctx1),
.data_in_ctx2(MEMC96_data_in_ctx2),
.data_out_ctx1(MEMC96_data_out_ctx1),
.data_out_ctx2(MEMC96_data_out_ctx2),
.write_mem_en_ctx1(MEMC96_write_mem_en_ctx1),
.mem_en_ctx1(MEMC96_mem_en_ctx1),.write_mem_en_ctx2(MEMC96_write_mem_en_ctx2),
.mem_en_ctx2(MEMC96_mem_en_ctx2));

defparam MEMC96.DATA_WIDTH = 32;
defparam MEMC96.ADDR_WIDTH = 6;
defparam MEMC96.STRIDE_WIDTH = 1;
wire MEMC97_valid_ctx1;
wire MEMC97_valid_ctx2;
wire [31:0] MEMC97_data_from_Core;
wire [31:0] MEMC97_data_to_Core;
wire [5:0] MEMC97_addr_out_ctx1;
wire MEMC97_write_en_ctx1;
wire MEMC97_write_mem_en_ctx1;
wire MEMC97_mem_en_ctx1;
wire [5:0] MEMC97_start_addr_ctx1;
wire [0:0] MEMC97_stride_ctx1;
wire [5:0] MEMC97_addr_out_ctx2;
wire MEMC97_write_en_ctx2;
wire MEMC97_write_mem_en_ctx2;
wire MEMC97_mem_en_ctx2;
wire [5:0] MEMC97_start_addr_ctx2;
wire [0:0] MEMC97_stride_ctx2;
wire [31:0] MEMC97_data_in_ctx1;
wire [31:0] MEMC97_data_in_ctx2;
wire [31:0] MEMC97_data_out_ctx1;
wire [31:0] MEMC97_data_out_ctx2;
wire [63:0] MEMC97_burst_count_ctx1;
wire [63:0] MEMC97_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC97(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC97_data_from_Core),
.data_to_Core(MEMC97_data_to_Core),
.valid_ctx1(MEMC97_valid_ctx1),
.addr_out_ctx1(MEMC97_addr_out_ctx1),
.write_en_ctx1(MEMC97_write_en_ctx1),
.start_addr_ctx1(MEMC97_start_addr_ctx1),
.stride_ctx1(MEMC97_stride_ctx1),
.burst_count_ctx1(MEMC97_burst_count_ctx1),
.valid_ctx2(MEMC97_valid_ctx2),
.addr_out_ctx2(MEMC97_addr_out_ctx2),
.write_en_ctx2(MEMC97_write_en_ctx2),
.start_addr_ctx2(MEMC97_start_addr_ctx2),
.stride_ctx2(MEMC97_stride_ctx2),
.burst_count_ctx2(MEMC97_burst_count_ctx2),
.data_in_ctx1(MEMC97_data_in_ctx1),
.data_in_ctx2(MEMC97_data_in_ctx2),
.data_out_ctx1(MEMC97_data_out_ctx1),
.data_out_ctx2(MEMC97_data_out_ctx2),
.write_mem_en_ctx1(MEMC97_write_mem_en_ctx1),
.mem_en_ctx1(MEMC97_mem_en_ctx1),.write_mem_en_ctx2(MEMC97_write_mem_en_ctx2),
.mem_en_ctx2(MEMC97_mem_en_ctx2));

defparam MEMC97.DATA_WIDTH = 32;
defparam MEMC97.ADDR_WIDTH = 6;
defparam MEMC97.STRIDE_WIDTH = 1;
wire MEMC98_valid_ctx1;
wire MEMC98_valid_ctx2;
wire [31:0] MEMC98_data_from_Core;
wire [31:0] MEMC98_data_to_Core;
wire [5:0] MEMC98_addr_out_ctx1;
wire MEMC98_write_en_ctx1;
wire MEMC98_write_mem_en_ctx1;
wire MEMC98_mem_en_ctx1;
wire [5:0] MEMC98_start_addr_ctx1;
wire [0:0] MEMC98_stride_ctx1;
wire [5:0] MEMC98_addr_out_ctx2;
wire MEMC98_write_en_ctx2;
wire MEMC98_write_mem_en_ctx2;
wire MEMC98_mem_en_ctx2;
wire [5:0] MEMC98_start_addr_ctx2;
wire [0:0] MEMC98_stride_ctx2;
wire [31:0] MEMC98_data_in_ctx1;
wire [31:0] MEMC98_data_in_ctx2;
wire [31:0] MEMC98_data_out_ctx1;
wire [31:0] MEMC98_data_out_ctx2;
wire [63:0] MEMC98_burst_count_ctx1;
wire [63:0] MEMC98_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC98(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC98_data_from_Core),
.data_to_Core(MEMC98_data_to_Core),
.valid_ctx1(MEMC98_valid_ctx1),
.addr_out_ctx1(MEMC98_addr_out_ctx1),
.write_en_ctx1(MEMC98_write_en_ctx1),
.start_addr_ctx1(MEMC98_start_addr_ctx1),
.stride_ctx1(MEMC98_stride_ctx1),
.burst_count_ctx1(MEMC98_burst_count_ctx1),
.valid_ctx2(MEMC98_valid_ctx2),
.addr_out_ctx2(MEMC98_addr_out_ctx2),
.write_en_ctx2(MEMC98_write_en_ctx2),
.start_addr_ctx2(MEMC98_start_addr_ctx2),
.stride_ctx2(MEMC98_stride_ctx2),
.burst_count_ctx2(MEMC98_burst_count_ctx2),
.data_in_ctx1(MEMC98_data_in_ctx1),
.data_in_ctx2(MEMC98_data_in_ctx2),
.data_out_ctx1(MEMC98_data_out_ctx1),
.data_out_ctx2(MEMC98_data_out_ctx2),
.write_mem_en_ctx1(MEMC98_write_mem_en_ctx1),
.mem_en_ctx1(MEMC98_mem_en_ctx1),.write_mem_en_ctx2(MEMC98_write_mem_en_ctx2),
.mem_en_ctx2(MEMC98_mem_en_ctx2));

defparam MEMC98.DATA_WIDTH = 32;
defparam MEMC98.ADDR_WIDTH = 6;
defparam MEMC98.STRIDE_WIDTH = 1;
wire MEMC99_valid_ctx1;
wire MEMC99_valid_ctx2;
wire [31:0] MEMC99_data_from_Core;
wire [31:0] MEMC99_data_to_Core;
wire [5:0] MEMC99_addr_out_ctx1;
wire MEMC99_write_en_ctx1;
wire MEMC99_write_mem_en_ctx1;
wire MEMC99_mem_en_ctx1;
wire [5:0] MEMC99_start_addr_ctx1;
wire [0:0] MEMC99_stride_ctx1;
wire [5:0] MEMC99_addr_out_ctx2;
wire MEMC99_write_en_ctx2;
wire MEMC99_write_mem_en_ctx2;
wire MEMC99_mem_en_ctx2;
wire [5:0] MEMC99_start_addr_ctx2;
wire [0:0] MEMC99_stride_ctx2;
wire [31:0] MEMC99_data_in_ctx1;
wire [31:0] MEMC99_data_in_ctx2;
wire [31:0] MEMC99_data_out_ctx1;
wire [31:0] MEMC99_data_out_ctx2;
wire [63:0] MEMC99_burst_count_ctx1;
wire [63:0] MEMC99_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC99(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC99_data_from_Core),
.data_to_Core(MEMC99_data_to_Core),
.valid_ctx1(MEMC99_valid_ctx1),
.addr_out_ctx1(MEMC99_addr_out_ctx1),
.write_en_ctx1(MEMC99_write_en_ctx1),
.start_addr_ctx1(MEMC99_start_addr_ctx1),
.stride_ctx1(MEMC99_stride_ctx1),
.burst_count_ctx1(MEMC99_burst_count_ctx1),
.valid_ctx2(MEMC99_valid_ctx2),
.addr_out_ctx2(MEMC99_addr_out_ctx2),
.write_en_ctx2(MEMC99_write_en_ctx2),
.start_addr_ctx2(MEMC99_start_addr_ctx2),
.stride_ctx2(MEMC99_stride_ctx2),
.burst_count_ctx2(MEMC99_burst_count_ctx2),
.data_in_ctx1(MEMC99_data_in_ctx1),
.data_in_ctx2(MEMC99_data_in_ctx2),
.data_out_ctx1(MEMC99_data_out_ctx1),
.data_out_ctx2(MEMC99_data_out_ctx2),
.write_mem_en_ctx1(MEMC99_write_mem_en_ctx1),
.mem_en_ctx1(MEMC99_mem_en_ctx1),.write_mem_en_ctx2(MEMC99_write_mem_en_ctx2),
.mem_en_ctx2(MEMC99_mem_en_ctx2));

defparam MEMC99.DATA_WIDTH = 32;
defparam MEMC99.ADDR_WIDTH = 6;
defparam MEMC99.STRIDE_WIDTH = 1;
wire MEMC100_valid_ctx1;
wire MEMC100_valid_ctx2;
wire [31:0] MEMC100_data_from_Core;
wire [31:0] MEMC100_data_to_Core;
wire [5:0] MEMC100_addr_out_ctx1;
wire MEMC100_write_en_ctx1;
wire MEMC100_write_mem_en_ctx1;
wire MEMC100_mem_en_ctx1;
wire [5:0] MEMC100_start_addr_ctx1;
wire [0:0] MEMC100_stride_ctx1;
wire [5:0] MEMC100_addr_out_ctx2;
wire MEMC100_write_en_ctx2;
wire MEMC100_write_mem_en_ctx2;
wire MEMC100_mem_en_ctx2;
wire [5:0] MEMC100_start_addr_ctx2;
wire [0:0] MEMC100_stride_ctx2;
wire [31:0] MEMC100_data_in_ctx1;
wire [31:0] MEMC100_data_in_ctx2;
wire [31:0] MEMC100_data_out_ctx1;
wire [31:0] MEMC100_data_out_ctx2;
wire [63:0] MEMC100_burst_count_ctx1;
wire [63:0] MEMC100_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC100(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC100_data_from_Core),
.data_to_Core(MEMC100_data_to_Core),
.valid_ctx1(MEMC100_valid_ctx1),
.addr_out_ctx1(MEMC100_addr_out_ctx1),
.write_en_ctx1(MEMC100_write_en_ctx1),
.start_addr_ctx1(MEMC100_start_addr_ctx1),
.stride_ctx1(MEMC100_stride_ctx1),
.burst_count_ctx1(MEMC100_burst_count_ctx1),
.valid_ctx2(MEMC100_valid_ctx2),
.addr_out_ctx2(MEMC100_addr_out_ctx2),
.write_en_ctx2(MEMC100_write_en_ctx2),
.start_addr_ctx2(MEMC100_start_addr_ctx2),
.stride_ctx2(MEMC100_stride_ctx2),
.burst_count_ctx2(MEMC100_burst_count_ctx2),
.data_in_ctx1(MEMC100_data_in_ctx1),
.data_in_ctx2(MEMC100_data_in_ctx2),
.data_out_ctx1(MEMC100_data_out_ctx1),
.data_out_ctx2(MEMC100_data_out_ctx2),
.write_mem_en_ctx1(MEMC100_write_mem_en_ctx1),
.mem_en_ctx1(MEMC100_mem_en_ctx1),.write_mem_en_ctx2(MEMC100_write_mem_en_ctx2),
.mem_en_ctx2(MEMC100_mem_en_ctx2));

defparam MEMC100.DATA_WIDTH = 32;
defparam MEMC100.ADDR_WIDTH = 6;
defparam MEMC100.STRIDE_WIDTH = 1;
wire MEMC101_valid_ctx1;
wire MEMC101_valid_ctx2;
wire [31:0] MEMC101_data_from_Core;
wire [31:0] MEMC101_data_to_Core;
wire [5:0] MEMC101_addr_out_ctx1;
wire MEMC101_write_en_ctx1;
wire MEMC101_write_mem_en_ctx1;
wire MEMC101_mem_en_ctx1;
wire [5:0] MEMC101_start_addr_ctx1;
wire [0:0] MEMC101_stride_ctx1;
wire [5:0] MEMC101_addr_out_ctx2;
wire MEMC101_write_en_ctx2;
wire MEMC101_write_mem_en_ctx2;
wire MEMC101_mem_en_ctx2;
wire [5:0] MEMC101_start_addr_ctx2;
wire [0:0] MEMC101_stride_ctx2;
wire [31:0] MEMC101_data_in_ctx1;
wire [31:0] MEMC101_data_in_ctx2;
wire [31:0] MEMC101_data_out_ctx1;
wire [31:0] MEMC101_data_out_ctx2;
wire [63:0] MEMC101_burst_count_ctx1;
wire [63:0] MEMC101_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC101(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC101_data_from_Core),
.data_to_Core(MEMC101_data_to_Core),
.valid_ctx1(MEMC101_valid_ctx1),
.addr_out_ctx1(MEMC101_addr_out_ctx1),
.write_en_ctx1(MEMC101_write_en_ctx1),
.start_addr_ctx1(MEMC101_start_addr_ctx1),
.stride_ctx1(MEMC101_stride_ctx1),
.burst_count_ctx1(MEMC101_burst_count_ctx1),
.valid_ctx2(MEMC101_valid_ctx2),
.addr_out_ctx2(MEMC101_addr_out_ctx2),
.write_en_ctx2(MEMC101_write_en_ctx2),
.start_addr_ctx2(MEMC101_start_addr_ctx2),
.stride_ctx2(MEMC101_stride_ctx2),
.burst_count_ctx2(MEMC101_burst_count_ctx2),
.data_in_ctx1(MEMC101_data_in_ctx1),
.data_in_ctx2(MEMC101_data_in_ctx2),
.data_out_ctx1(MEMC101_data_out_ctx1),
.data_out_ctx2(MEMC101_data_out_ctx2),
.write_mem_en_ctx1(MEMC101_write_mem_en_ctx1),
.mem_en_ctx1(MEMC101_mem_en_ctx1),.write_mem_en_ctx2(MEMC101_write_mem_en_ctx2),
.mem_en_ctx2(MEMC101_mem_en_ctx2));

defparam MEMC101.DATA_WIDTH = 32;
defparam MEMC101.ADDR_WIDTH = 6;
defparam MEMC101.STRIDE_WIDTH = 1;
wire MEMC102_valid_ctx1;
wire MEMC102_valid_ctx2;
wire [31:0] MEMC102_data_from_Core;
wire [31:0] MEMC102_data_to_Core;
wire [5:0] MEMC102_addr_out_ctx1;
wire MEMC102_write_en_ctx1;
wire MEMC102_write_mem_en_ctx1;
wire MEMC102_mem_en_ctx1;
wire [5:0] MEMC102_start_addr_ctx1;
wire [0:0] MEMC102_stride_ctx1;
wire [5:0] MEMC102_addr_out_ctx2;
wire MEMC102_write_en_ctx2;
wire MEMC102_write_mem_en_ctx2;
wire MEMC102_mem_en_ctx2;
wire [5:0] MEMC102_start_addr_ctx2;
wire [0:0] MEMC102_stride_ctx2;
wire [31:0] MEMC102_data_in_ctx1;
wire [31:0] MEMC102_data_in_ctx2;
wire [31:0] MEMC102_data_out_ctx1;
wire [31:0] MEMC102_data_out_ctx2;
wire [63:0] MEMC102_burst_count_ctx1;
wire [63:0] MEMC102_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC102(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC102_data_from_Core),
.data_to_Core(MEMC102_data_to_Core),
.valid_ctx1(MEMC102_valid_ctx1),
.addr_out_ctx1(MEMC102_addr_out_ctx1),
.write_en_ctx1(MEMC102_write_en_ctx1),
.start_addr_ctx1(MEMC102_start_addr_ctx1),
.stride_ctx1(MEMC102_stride_ctx1),
.burst_count_ctx1(MEMC102_burst_count_ctx1),
.valid_ctx2(MEMC102_valid_ctx2),
.addr_out_ctx2(MEMC102_addr_out_ctx2),
.write_en_ctx2(MEMC102_write_en_ctx2),
.start_addr_ctx2(MEMC102_start_addr_ctx2),
.stride_ctx2(MEMC102_stride_ctx2),
.burst_count_ctx2(MEMC102_burst_count_ctx2),
.data_in_ctx1(MEMC102_data_in_ctx1),
.data_in_ctx2(MEMC102_data_in_ctx2),
.data_out_ctx1(MEMC102_data_out_ctx1),
.data_out_ctx2(MEMC102_data_out_ctx2),
.write_mem_en_ctx1(MEMC102_write_mem_en_ctx1),
.mem_en_ctx1(MEMC102_mem_en_ctx1),.write_mem_en_ctx2(MEMC102_write_mem_en_ctx2),
.mem_en_ctx2(MEMC102_mem_en_ctx2));

defparam MEMC102.DATA_WIDTH = 32;
defparam MEMC102.ADDR_WIDTH = 6;
defparam MEMC102.STRIDE_WIDTH = 1;
wire MEMC103_valid_ctx1;
wire MEMC103_valid_ctx2;
wire [31:0] MEMC103_data_from_Core;
wire [31:0] MEMC103_data_to_Core;
wire [5:0] MEMC103_addr_out_ctx1;
wire MEMC103_write_en_ctx1;
wire MEMC103_write_mem_en_ctx1;
wire MEMC103_mem_en_ctx1;
wire [5:0] MEMC103_start_addr_ctx1;
wire [0:0] MEMC103_stride_ctx1;
wire [5:0] MEMC103_addr_out_ctx2;
wire MEMC103_write_en_ctx2;
wire MEMC103_write_mem_en_ctx2;
wire MEMC103_mem_en_ctx2;
wire [5:0] MEMC103_start_addr_ctx2;
wire [0:0] MEMC103_stride_ctx2;
wire [31:0] MEMC103_data_in_ctx1;
wire [31:0] MEMC103_data_in_ctx2;
wire [31:0] MEMC103_data_out_ctx1;
wire [31:0] MEMC103_data_out_ctx2;
wire [63:0] MEMC103_burst_count_ctx1;
wire [63:0] MEMC103_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC103(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC103_data_from_Core),
.data_to_Core(MEMC103_data_to_Core),
.valid_ctx1(MEMC103_valid_ctx1),
.addr_out_ctx1(MEMC103_addr_out_ctx1),
.write_en_ctx1(MEMC103_write_en_ctx1),
.start_addr_ctx1(MEMC103_start_addr_ctx1),
.stride_ctx1(MEMC103_stride_ctx1),
.burst_count_ctx1(MEMC103_burst_count_ctx1),
.valid_ctx2(MEMC103_valid_ctx2),
.addr_out_ctx2(MEMC103_addr_out_ctx2),
.write_en_ctx2(MEMC103_write_en_ctx2),
.start_addr_ctx2(MEMC103_start_addr_ctx2),
.stride_ctx2(MEMC103_stride_ctx2),
.burst_count_ctx2(MEMC103_burst_count_ctx2),
.data_in_ctx1(MEMC103_data_in_ctx1),
.data_in_ctx2(MEMC103_data_in_ctx2),
.data_out_ctx1(MEMC103_data_out_ctx1),
.data_out_ctx2(MEMC103_data_out_ctx2),
.write_mem_en_ctx1(MEMC103_write_mem_en_ctx1),
.mem_en_ctx1(MEMC103_mem_en_ctx1),.write_mem_en_ctx2(MEMC103_write_mem_en_ctx2),
.mem_en_ctx2(MEMC103_mem_en_ctx2));

defparam MEMC103.DATA_WIDTH = 32;
defparam MEMC103.ADDR_WIDTH = 6;
defparam MEMC103.STRIDE_WIDTH = 1;
wire MEMC104_valid_ctx1;
wire MEMC104_valid_ctx2;
wire [31:0] MEMC104_data_from_Core;
wire [31:0] MEMC104_data_to_Core;
wire [5:0] MEMC104_addr_out_ctx1;
wire MEMC104_write_en_ctx1;
wire MEMC104_write_mem_en_ctx1;
wire MEMC104_mem_en_ctx1;
wire [5:0] MEMC104_start_addr_ctx1;
wire [0:0] MEMC104_stride_ctx1;
wire [5:0] MEMC104_addr_out_ctx2;
wire MEMC104_write_en_ctx2;
wire MEMC104_write_mem_en_ctx2;
wire MEMC104_mem_en_ctx2;
wire [5:0] MEMC104_start_addr_ctx2;
wire [0:0] MEMC104_stride_ctx2;
wire [31:0] MEMC104_data_in_ctx1;
wire [31:0] MEMC104_data_in_ctx2;
wire [31:0] MEMC104_data_out_ctx1;
wire [31:0] MEMC104_data_out_ctx2;
wire [63:0] MEMC104_burst_count_ctx1;
wire [63:0] MEMC104_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC104(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC104_data_from_Core),
.data_to_Core(MEMC104_data_to_Core),
.valid_ctx1(MEMC104_valid_ctx1),
.addr_out_ctx1(MEMC104_addr_out_ctx1),
.write_en_ctx1(MEMC104_write_en_ctx1),
.start_addr_ctx1(MEMC104_start_addr_ctx1),
.stride_ctx1(MEMC104_stride_ctx1),
.burst_count_ctx1(MEMC104_burst_count_ctx1),
.valid_ctx2(MEMC104_valid_ctx2),
.addr_out_ctx2(MEMC104_addr_out_ctx2),
.write_en_ctx2(MEMC104_write_en_ctx2),
.start_addr_ctx2(MEMC104_start_addr_ctx2),
.stride_ctx2(MEMC104_stride_ctx2),
.burst_count_ctx2(MEMC104_burst_count_ctx2),
.data_in_ctx1(MEMC104_data_in_ctx1),
.data_in_ctx2(MEMC104_data_in_ctx2),
.data_out_ctx1(MEMC104_data_out_ctx1),
.data_out_ctx2(MEMC104_data_out_ctx2),
.write_mem_en_ctx1(MEMC104_write_mem_en_ctx1),
.mem_en_ctx1(MEMC104_mem_en_ctx1),.write_mem_en_ctx2(MEMC104_write_mem_en_ctx2),
.mem_en_ctx2(MEMC104_mem_en_ctx2));

defparam MEMC104.DATA_WIDTH = 32;
defparam MEMC104.ADDR_WIDTH = 6;
defparam MEMC104.STRIDE_WIDTH = 1;
wire MEMC105_valid_ctx1;
wire MEMC105_valid_ctx2;
wire [31:0] MEMC105_data_from_Core;
wire [31:0] MEMC105_data_to_Core;
wire [5:0] MEMC105_addr_out_ctx1;
wire MEMC105_write_en_ctx1;
wire MEMC105_write_mem_en_ctx1;
wire MEMC105_mem_en_ctx1;
wire [5:0] MEMC105_start_addr_ctx1;
wire [0:0] MEMC105_stride_ctx1;
wire [5:0] MEMC105_addr_out_ctx2;
wire MEMC105_write_en_ctx2;
wire MEMC105_write_mem_en_ctx2;
wire MEMC105_mem_en_ctx2;
wire [5:0] MEMC105_start_addr_ctx2;
wire [0:0] MEMC105_stride_ctx2;
wire [31:0] MEMC105_data_in_ctx1;
wire [31:0] MEMC105_data_in_ctx2;
wire [31:0] MEMC105_data_out_ctx1;
wire [31:0] MEMC105_data_out_ctx2;
wire [63:0] MEMC105_burst_count_ctx1;
wire [63:0] MEMC105_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC105(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC105_data_from_Core),
.data_to_Core(MEMC105_data_to_Core),
.valid_ctx1(MEMC105_valid_ctx1),
.addr_out_ctx1(MEMC105_addr_out_ctx1),
.write_en_ctx1(MEMC105_write_en_ctx1),
.start_addr_ctx1(MEMC105_start_addr_ctx1),
.stride_ctx1(MEMC105_stride_ctx1),
.burst_count_ctx1(MEMC105_burst_count_ctx1),
.valid_ctx2(MEMC105_valid_ctx2),
.addr_out_ctx2(MEMC105_addr_out_ctx2),
.write_en_ctx2(MEMC105_write_en_ctx2),
.start_addr_ctx2(MEMC105_start_addr_ctx2),
.stride_ctx2(MEMC105_stride_ctx2),
.burst_count_ctx2(MEMC105_burst_count_ctx2),
.data_in_ctx1(MEMC105_data_in_ctx1),
.data_in_ctx2(MEMC105_data_in_ctx2),
.data_out_ctx1(MEMC105_data_out_ctx1),
.data_out_ctx2(MEMC105_data_out_ctx2),
.write_mem_en_ctx1(MEMC105_write_mem_en_ctx1),
.mem_en_ctx1(MEMC105_mem_en_ctx1),.write_mem_en_ctx2(MEMC105_write_mem_en_ctx2),
.mem_en_ctx2(MEMC105_mem_en_ctx2));

defparam MEMC105.DATA_WIDTH = 32;
defparam MEMC105.ADDR_WIDTH = 6;
defparam MEMC105.STRIDE_WIDTH = 1;
wire MEMC106_valid_ctx1;
wire MEMC106_valid_ctx2;
wire [31:0] MEMC106_data_from_Core;
wire [31:0] MEMC106_data_to_Core;
wire [5:0] MEMC106_addr_out_ctx1;
wire MEMC106_write_en_ctx1;
wire MEMC106_write_mem_en_ctx1;
wire MEMC106_mem_en_ctx1;
wire [5:0] MEMC106_start_addr_ctx1;
wire [0:0] MEMC106_stride_ctx1;
wire [5:0] MEMC106_addr_out_ctx2;
wire MEMC106_write_en_ctx2;
wire MEMC106_write_mem_en_ctx2;
wire MEMC106_mem_en_ctx2;
wire [5:0] MEMC106_start_addr_ctx2;
wire [0:0] MEMC106_stride_ctx2;
wire [31:0] MEMC106_data_in_ctx1;
wire [31:0] MEMC106_data_in_ctx2;
wire [31:0] MEMC106_data_out_ctx1;
wire [31:0] MEMC106_data_out_ctx2;
wire [63:0] MEMC106_burst_count_ctx1;
wire [63:0] MEMC106_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC106(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC106_data_from_Core),
.data_to_Core(MEMC106_data_to_Core),
.valid_ctx1(MEMC106_valid_ctx1),
.addr_out_ctx1(MEMC106_addr_out_ctx1),
.write_en_ctx1(MEMC106_write_en_ctx1),
.start_addr_ctx1(MEMC106_start_addr_ctx1),
.stride_ctx1(MEMC106_stride_ctx1),
.burst_count_ctx1(MEMC106_burst_count_ctx1),
.valid_ctx2(MEMC106_valid_ctx2),
.addr_out_ctx2(MEMC106_addr_out_ctx2),
.write_en_ctx2(MEMC106_write_en_ctx2),
.start_addr_ctx2(MEMC106_start_addr_ctx2),
.stride_ctx2(MEMC106_stride_ctx2),
.burst_count_ctx2(MEMC106_burst_count_ctx2),
.data_in_ctx1(MEMC106_data_in_ctx1),
.data_in_ctx2(MEMC106_data_in_ctx2),
.data_out_ctx1(MEMC106_data_out_ctx1),
.data_out_ctx2(MEMC106_data_out_ctx2),
.write_mem_en_ctx1(MEMC106_write_mem_en_ctx1),
.mem_en_ctx1(MEMC106_mem_en_ctx1),.write_mem_en_ctx2(MEMC106_write_mem_en_ctx2),
.mem_en_ctx2(MEMC106_mem_en_ctx2));

defparam MEMC106.DATA_WIDTH = 32;
defparam MEMC106.ADDR_WIDTH = 6;
defparam MEMC106.STRIDE_WIDTH = 1;
wire MEMC107_valid_ctx1;
wire MEMC107_valid_ctx2;
wire [31:0] MEMC107_data_from_Core;
wire [31:0] MEMC107_data_to_Core;
wire [5:0] MEMC107_addr_out_ctx1;
wire MEMC107_write_en_ctx1;
wire MEMC107_write_mem_en_ctx1;
wire MEMC107_mem_en_ctx1;
wire [5:0] MEMC107_start_addr_ctx1;
wire [0:0] MEMC107_stride_ctx1;
wire [5:0] MEMC107_addr_out_ctx2;
wire MEMC107_write_en_ctx2;
wire MEMC107_write_mem_en_ctx2;
wire MEMC107_mem_en_ctx2;
wire [5:0] MEMC107_start_addr_ctx2;
wire [0:0] MEMC107_stride_ctx2;
wire [31:0] MEMC107_data_in_ctx1;
wire [31:0] MEMC107_data_in_ctx2;
wire [31:0] MEMC107_data_out_ctx1;
wire [31:0] MEMC107_data_out_ctx2;
wire [63:0] MEMC107_burst_count_ctx1;
wire [63:0] MEMC107_burst_count_ctx2;
CADA_TDP_MemControlBurst MEMC107(
.clk(clk),
.rst(rst),
.data_from_Core(MEMC107_data_from_Core),
.data_to_Core(MEMC107_data_to_Core),
.valid_ctx1(MEMC107_valid_ctx1),
.addr_out_ctx1(MEMC107_addr_out_ctx1),
.write_en_ctx1(MEMC107_write_en_ctx1),
.start_addr_ctx1(MEMC107_start_addr_ctx1),
.stride_ctx1(MEMC107_stride_ctx1),
.burst_count_ctx1(MEMC107_burst_count_ctx1),
.valid_ctx2(MEMC107_valid_ctx2),
.addr_out_ctx2(MEMC107_addr_out_ctx2),
.write_en_ctx2(MEMC107_write_en_ctx2),
.start_addr_ctx2(MEMC107_start_addr_ctx2),
.stride_ctx2(MEMC107_stride_ctx2),
.burst_count_ctx2(MEMC107_burst_count_ctx2),
.data_in_ctx1(MEMC107_data_in_ctx1),
.data_in_ctx2(MEMC107_data_in_ctx2),
.data_out_ctx1(MEMC107_data_out_ctx1),
.data_out_ctx2(MEMC107_data_out_ctx2),
.write_mem_en_ctx1(MEMC107_write_mem_en_ctx1),
.mem_en_ctx1(MEMC107_mem_en_ctx1),.write_mem_en_ctx2(MEMC107_write_mem_en_ctx2),
.mem_en_ctx2(MEMC107_mem_en_ctx2));

defparam MEMC107.DATA_WIDTH = 32;
defparam MEMC107.ADDR_WIDTH = 6;
defparam MEMC107.STRIDE_WIDTH = 1;
wire IMEMC_valid_ctx1;
wire IMEMC_valid_ctx2;
wire [38:0] IMEMC_data_to_Core;
wire [38:0] IMEMC_data_from_Core;
wire [4:0] IMEMC_addr_out_ctx1;
wire IMEMC_write_en_ctx1;
wire IMEMC_mem_en_ctx1;
wire IMEMC_write_mem_en_ctx1;
wire [4:0] IMEMC_start_addr_ctx1;
wire [0:0] IMEMC_stride_ctx1;
wire [38:0] IMEMC_data_in_ctx1;
wire [38:0] IMEMC_data_in_ctx2;
wire [38:0] IMEMC_data_out_ctx1;
wire [38:0] IMEMC_data_out_ctx2;
wire [4:0] IMEMC_addr_out_ctx2;
wire IMEMC_write_en_ctx2;
wire IMEMC_mem_en_ctx2;
wire IMEMC_write_mem_en_ctx2;
wire [4:0] IMEMC_start_addr_ctx2;
wire [0:0] IMEMC_stride_ctx2;
wire [199:0] IMEMC_burst_count_ctx1;
wire [199:0] IMEMC_burst_count_ctx2;
CADA_TDP_MemControlBurst IMEMC(
.clk(clk),
.rst(rst),
.data_from_Core(IMEMC_data_from_Core),
.data_to_Core(IMEMC_data_to_Core),
.valid_ctx1(IMEMC_valid_ctx1),
.addr_out_ctx1(IMEMC_addr_out_ctx1),
.write_en_ctx1(IMEMC_write_en_ctx1),
.start_addr_ctx1(IMEMC_start_addr_ctx1),
.stride_ctx1(IMEMC_stride_ctx1),
.burst_count_ctx1(IMEMC_burst_count_ctx1),
.valid_ctx2(IMEMC_valid_ctx2),
.addr_out_ctx2(IMEMC_addr_out_ctx2),
.write_en_ctx2(IMEMC_write_en_ctx2),
.start_addr_ctx2(IMEMC_start_addr_ctx2),
.stride_ctx2(IMEMC_stride_ctx2),
.burst_count_ctx2(IMEMC_burst_count_ctx2),
.data_in_ctx1(IMEMC_data_in_ctx1),
.data_in_ctx2(IMEMC_data_in_ctx2),
.data_out_ctx1(IMEMC_data_out_ctx1),
.data_out_ctx2(IMEMC_data_out_ctx2),
.write_mem_en_ctx1(IMEMC_write_mem_en_ctx1),
.mem_en_ctx1(IMEMC_mem_en_ctx1),.write_mem_en_ctx2(IMEMC_write_mem_en_ctx2),
.mem_en_ctx2(IMEMC_mem_en_ctx2));

defparam IMEMC.DATA_WIDTH = 39;
defparam IMEMC.ADDR_WIDTH = 5;
defparam IMEMC.STRIDE_WIDTH = 1;
assign gControlInW = IOConfig[125:0];

assign mOutConfigW = IOConfig[557:126];

assign controlInW = IMEMC_data_to_Core[35:0]; 

assign configInW = IMEMC_data_to_Core[38:36]; 

wire [31:0] MEMOCMux0_inw1;
wire [31:0] MEMOCMux0_inw2;
wire [31:0] MEMOCMux0_inw3;
wire [31:0] MEMOCMux0_inw4;
wire [31:0] MEMOCMux0_inw5;
wire [31:0] MEMOCMux0_inw6;
wire [31:0] MEMOCMux0_inw7;
wire [31:0] MEMOCMux0_inw8;
wire [31:0] MEMOCMux0_inw9;
wire [31:0] MEMOCMux0_inw10;
wire [31:0] MEMOCMux0_outw1;
wire [3:0] MEMOCMux0_selw;
HA_10IM MEMOCMux0 (
.DataIn_1(MEMOCMux0_inw1),
.DataIn_2(MEMOCMux0_inw2),
.DataIn_3(MEMOCMux0_inw3),
.DataIn_4(MEMOCMux0_inw4),
.DataIn_5(MEMOCMux0_inw5),
.DataIn_6(MEMOCMux0_inw6),
.DataIn_7(MEMOCMux0_inw7),
.DataIn_8(MEMOCMux0_inw8),
.DataIn_9(MEMOCMux0_inw9),
.DataIn_10(MEMOCMux0_inw10),
.DataOut_1(MEMOCMux0_outw1),
.sel(MEMOCMux0_selw));
defparam MEMOCMux0.Mux_BW = 32;
assign MEMC0_data_from_Core = MEMOCMux0_outw1;
assign MEMOCMux0_inw1 = dataOutW[31:0]; 
assign MEMOCMux0_inw2 = dataOutW[63:32]; 
assign MEMOCMux0_inw3 = dataOutW[95:64]; 
assign MEMOCMux0_inw4 = dataOutW[127:96]; 
assign MEMOCMux0_inw5 = dataOutW[159:128]; 
assign MEMOCMux0_inw6 = dataOutW[191:160]; 
assign MEMOCMux0_inw7 = dataOutW[223:192]; 
assign MEMOCMux0_inw8 = dataOutW[255:224]; 
assign MEMOCMux0_inw9 = dataOutW[287:256]; 
assign MEMOCMux0_inw10 = globalDataIn[31:0]; 
assign MEMOCMux0_selw = mOutConfigW[3:0]; 
assign MEMC0_data_out_ctx2 = mDataFromMem[31:0]; 
assign mDataToMem[31:0] = MEMC0_data_in_ctx1; 
assign globalDataOut[31:0] = MEMC0_data_to_Core; 
assign MEMC0_valid_ctx1 = valid1[0:0]; 
assign MEMC0_write_en_ctx1 = WEn1[0:0]; 
assign MEMC0_stride_ctx1 = stride1[0:0]; 
assign MEMC0_start_addr_ctx1 = startAddr1[5:0]; 
assign MEMC0_burst_count_ctx1 = count1[6:0]; 
assign mAddr1[5:0] = MEMC0_addr_out_ctx1; 
assign mEn1[0:0] = MEMC0_mem_en_ctx1; 
assign mWEn1[0:0] = MEMC0_write_mem_en_ctx1; 
assign MEMC0_valid_ctx2 = valid2[0:0]; 
assign MEMC0_write_en_ctx2 = WEn2[0:0]; 
assign MEMC0_stride_ctx2 = stride2[0:0]; 
assign MEMC0_start_addr_ctx2 = startAddr2[5:0]; 
assign mAddr2[5:0] = MEMC0_addr_out_ctx2; 
assign MEMC0_burst_count_ctx2 = count2[6:0]; 
assign mEn2[0:0] = MEMC0_mem_en_ctx2; 
assign mWEn2[0:0] = MEMC0_write_mem_en_ctx2; 
wire [31:0] MEMOCMux1_inw1;
wire [31:0] MEMOCMux1_inw2;
wire [31:0] MEMOCMux1_inw3;
wire [31:0] MEMOCMux1_inw4;
wire [31:0] MEMOCMux1_inw5;
wire [31:0] MEMOCMux1_inw6;
wire [31:0] MEMOCMux1_inw7;
wire [31:0] MEMOCMux1_inw8;
wire [31:0] MEMOCMux1_inw9;
wire [31:0] MEMOCMux1_inw10;
wire [31:0] MEMOCMux1_outw1;
wire [3:0] MEMOCMux1_selw;
HA_10IM MEMOCMux1 (
.DataIn_1(MEMOCMux1_inw1),
.DataIn_2(MEMOCMux1_inw2),
.DataIn_3(MEMOCMux1_inw3),
.DataIn_4(MEMOCMux1_inw4),
.DataIn_5(MEMOCMux1_inw5),
.DataIn_6(MEMOCMux1_inw6),
.DataIn_7(MEMOCMux1_inw7),
.DataIn_8(MEMOCMux1_inw8),
.DataIn_9(MEMOCMux1_inw9),
.DataIn_10(MEMOCMux1_inw10),
.DataOut_1(MEMOCMux1_outw1),
.sel(MEMOCMux1_selw));
defparam MEMOCMux1.Mux_BW = 32;
assign MEMC1_data_from_Core = MEMOCMux1_outw1;
assign MEMOCMux1_inw1 = dataOutW[31:0]; 
assign MEMOCMux1_inw2 = dataOutW[63:32]; 
assign MEMOCMux1_inw3 = dataOutW[95:64]; 
assign MEMOCMux1_inw4 = dataOutW[127:96]; 
assign MEMOCMux1_inw5 = dataOutW[159:128]; 
assign MEMOCMux1_inw6 = dataOutW[191:160]; 
assign MEMOCMux1_inw7 = dataOutW[223:192]; 
assign MEMOCMux1_inw8 = dataOutW[255:224]; 
assign MEMOCMux1_inw9 = dataOutW[287:256]; 
assign MEMOCMux1_inw10 = globalDataIn[63:32]; 
assign MEMOCMux1_selw = mOutConfigW[7:4]; 
assign MEMC1_data_out_ctx2 = mDataFromMem[63:32]; 
assign mDataToMem[63:32] = MEMC1_data_in_ctx1; 
assign globalDataOut[63:32] = MEMC1_data_to_Core; 
assign MEMC1_valid_ctx1 = valid1[1:1]; 
assign MEMC1_write_en_ctx1 = WEn1[1:1]; 
assign MEMC1_stride_ctx1 = stride1[1:1]; 
assign MEMC1_start_addr_ctx1 = startAddr1[11:6]; 
assign MEMC1_burst_count_ctx1 = count1[13:7]; 
assign mAddr1[11:6] = MEMC1_addr_out_ctx1; 
assign mEn1[1:1] = MEMC1_mem_en_ctx1; 
assign mWEn1[1:1] = MEMC1_write_mem_en_ctx1; 
assign MEMC1_valid_ctx2 = valid2[1:1]; 
assign MEMC1_write_en_ctx2 = WEn2[1:1]; 
assign MEMC1_stride_ctx2 = stride2[1:1]; 
assign MEMC1_start_addr_ctx2 = startAddr2[11:6]; 
assign mAddr2[11:6] = MEMC1_addr_out_ctx2; 
assign MEMC1_burst_count_ctx2 = count2[13:7]; 
assign mEn2[1:1] = MEMC1_mem_en_ctx2; 
assign mWEn2[1:1] = MEMC1_write_mem_en_ctx2; 
wire [31:0] MEMOCMux2_inw1;
wire [31:0] MEMOCMux2_inw2;
wire [31:0] MEMOCMux2_inw3;
wire [31:0] MEMOCMux2_inw4;
wire [31:0] MEMOCMux2_inw5;
wire [31:0] MEMOCMux2_inw6;
wire [31:0] MEMOCMux2_inw7;
wire [31:0] MEMOCMux2_inw8;
wire [31:0] MEMOCMux2_inw9;
wire [31:0] MEMOCMux2_inw10;
wire [31:0] MEMOCMux2_outw1;
wire [3:0] MEMOCMux2_selw;
HA_10IM MEMOCMux2 (
.DataIn_1(MEMOCMux2_inw1),
.DataIn_2(MEMOCMux2_inw2),
.DataIn_3(MEMOCMux2_inw3),
.DataIn_4(MEMOCMux2_inw4),
.DataIn_5(MEMOCMux2_inw5),
.DataIn_6(MEMOCMux2_inw6),
.DataIn_7(MEMOCMux2_inw7),
.DataIn_8(MEMOCMux2_inw8),
.DataIn_9(MEMOCMux2_inw9),
.DataIn_10(MEMOCMux2_inw10),
.DataOut_1(MEMOCMux2_outw1),
.sel(MEMOCMux2_selw));
defparam MEMOCMux2.Mux_BW = 32;
assign MEMC2_data_from_Core = MEMOCMux2_outw1;
assign MEMOCMux2_inw1 = dataOutW[31:0]; 
assign MEMOCMux2_inw2 = dataOutW[63:32]; 
assign MEMOCMux2_inw3 = dataOutW[95:64]; 
assign MEMOCMux2_inw4 = dataOutW[127:96]; 
assign MEMOCMux2_inw5 = dataOutW[159:128]; 
assign MEMOCMux2_inw6 = dataOutW[191:160]; 
assign MEMOCMux2_inw7 = dataOutW[223:192]; 
assign MEMOCMux2_inw8 = dataOutW[255:224]; 
assign MEMOCMux2_inw9 = dataOutW[287:256]; 
assign MEMOCMux2_inw10 = globalDataIn[95:64]; 
assign MEMOCMux2_selw = mOutConfigW[11:8]; 
assign MEMC2_data_out_ctx2 = mDataFromMem[95:64]; 
assign mDataToMem[95:64] = MEMC2_data_in_ctx1; 
assign globalDataOut[95:64] = MEMC2_data_to_Core; 
assign MEMC2_valid_ctx1 = valid1[2:2]; 
assign MEMC2_write_en_ctx1 = WEn1[2:2]; 
assign MEMC2_stride_ctx1 = stride1[2:2]; 
assign MEMC2_start_addr_ctx1 = startAddr1[17:12]; 
assign MEMC2_burst_count_ctx1 = count1[20:14]; 
assign mAddr1[17:12] = MEMC2_addr_out_ctx1; 
assign mEn1[2:2] = MEMC2_mem_en_ctx1; 
assign mWEn1[2:2] = MEMC2_write_mem_en_ctx1; 
assign MEMC2_valid_ctx2 = valid2[2:2]; 
assign MEMC2_write_en_ctx2 = WEn2[2:2]; 
assign MEMC2_stride_ctx2 = stride2[2:2]; 
assign MEMC2_start_addr_ctx2 = startAddr2[17:12]; 
assign mAddr2[17:12] = MEMC2_addr_out_ctx2; 
assign MEMC2_burst_count_ctx2 = count2[20:14]; 
assign mEn2[2:2] = MEMC2_mem_en_ctx2; 
assign mWEn2[2:2] = MEMC2_write_mem_en_ctx2; 
wire [31:0] MEMOCMux3_inw1;
wire [31:0] MEMOCMux3_inw2;
wire [31:0] MEMOCMux3_inw3;
wire [31:0] MEMOCMux3_inw4;
wire [31:0] MEMOCMux3_inw5;
wire [31:0] MEMOCMux3_inw6;
wire [31:0] MEMOCMux3_inw7;
wire [31:0] MEMOCMux3_inw8;
wire [31:0] MEMOCMux3_inw9;
wire [31:0] MEMOCMux3_inw10;
wire [31:0] MEMOCMux3_outw1;
wire [3:0] MEMOCMux3_selw;
HA_10IM MEMOCMux3 (
.DataIn_1(MEMOCMux3_inw1),
.DataIn_2(MEMOCMux3_inw2),
.DataIn_3(MEMOCMux3_inw3),
.DataIn_4(MEMOCMux3_inw4),
.DataIn_5(MEMOCMux3_inw5),
.DataIn_6(MEMOCMux3_inw6),
.DataIn_7(MEMOCMux3_inw7),
.DataIn_8(MEMOCMux3_inw8),
.DataIn_9(MEMOCMux3_inw9),
.DataIn_10(MEMOCMux3_inw10),
.DataOut_1(MEMOCMux3_outw1),
.sel(MEMOCMux3_selw));
defparam MEMOCMux3.Mux_BW = 32;
assign MEMC3_data_from_Core = MEMOCMux3_outw1;
assign MEMOCMux3_inw1 = dataOutW[31:0]; 
assign MEMOCMux3_inw2 = dataOutW[63:32]; 
assign MEMOCMux3_inw3 = dataOutW[95:64]; 
assign MEMOCMux3_inw4 = dataOutW[127:96]; 
assign MEMOCMux3_inw5 = dataOutW[159:128]; 
assign MEMOCMux3_inw6 = dataOutW[191:160]; 
assign MEMOCMux3_inw7 = dataOutW[223:192]; 
assign MEMOCMux3_inw8 = dataOutW[255:224]; 
assign MEMOCMux3_inw9 = dataOutW[287:256]; 
assign MEMOCMux3_inw10 = globalDataIn[127:96]; 
assign MEMOCMux3_selw = mOutConfigW[15:12]; 
assign MEMC3_data_out_ctx2 = mDataFromMem[127:96]; 
assign mDataToMem[127:96] = MEMC3_data_in_ctx1; 
assign globalDataOut[127:96] = MEMC3_data_to_Core; 
assign MEMC3_valid_ctx1 = valid1[3:3]; 
assign MEMC3_write_en_ctx1 = WEn1[3:3]; 
assign MEMC3_stride_ctx1 = stride1[3:3]; 
assign MEMC3_start_addr_ctx1 = startAddr1[23:18]; 
assign MEMC3_burst_count_ctx1 = count1[27:21]; 
assign mAddr1[23:18] = MEMC3_addr_out_ctx1; 
assign mEn1[3:3] = MEMC3_mem_en_ctx1; 
assign mWEn1[3:3] = MEMC3_write_mem_en_ctx1; 
assign MEMC3_valid_ctx2 = valid2[3:3]; 
assign MEMC3_write_en_ctx2 = WEn2[3:3]; 
assign MEMC3_stride_ctx2 = stride2[3:3]; 
assign MEMC3_start_addr_ctx2 = startAddr2[23:18]; 
assign mAddr2[23:18] = MEMC3_addr_out_ctx2; 
assign MEMC3_burst_count_ctx2 = count2[27:21]; 
assign mEn2[3:3] = MEMC3_mem_en_ctx2; 
assign mWEn2[3:3] = MEMC3_write_mem_en_ctx2; 
wire [31:0] MEMOCMux4_inw1;
wire [31:0] MEMOCMux4_inw2;
wire [31:0] MEMOCMux4_inw3;
wire [31:0] MEMOCMux4_inw4;
wire [31:0] MEMOCMux4_inw5;
wire [31:0] MEMOCMux4_inw6;
wire [31:0] MEMOCMux4_inw7;
wire [31:0] MEMOCMux4_inw8;
wire [31:0] MEMOCMux4_inw9;
wire [31:0] MEMOCMux4_inw10;
wire [31:0] MEMOCMux4_outw1;
wire [3:0] MEMOCMux4_selw;
HA_10IM MEMOCMux4 (
.DataIn_1(MEMOCMux4_inw1),
.DataIn_2(MEMOCMux4_inw2),
.DataIn_3(MEMOCMux4_inw3),
.DataIn_4(MEMOCMux4_inw4),
.DataIn_5(MEMOCMux4_inw5),
.DataIn_6(MEMOCMux4_inw6),
.DataIn_7(MEMOCMux4_inw7),
.DataIn_8(MEMOCMux4_inw8),
.DataIn_9(MEMOCMux4_inw9),
.DataIn_10(MEMOCMux4_inw10),
.DataOut_1(MEMOCMux4_outw1),
.sel(MEMOCMux4_selw));
defparam MEMOCMux4.Mux_BW = 32;
assign MEMC4_data_from_Core = MEMOCMux4_outw1;
assign MEMOCMux4_inw1 = dataOutW[31:0]; 
assign MEMOCMux4_inw2 = dataOutW[63:32]; 
assign MEMOCMux4_inw3 = dataOutW[95:64]; 
assign MEMOCMux4_inw4 = dataOutW[127:96]; 
assign MEMOCMux4_inw5 = dataOutW[159:128]; 
assign MEMOCMux4_inw6 = dataOutW[191:160]; 
assign MEMOCMux4_inw7 = dataOutW[223:192]; 
assign MEMOCMux4_inw8 = dataOutW[255:224]; 
assign MEMOCMux4_inw9 = dataOutW[287:256]; 
assign MEMOCMux4_inw10 = globalDataIn[159:128]; 
assign MEMOCMux4_selw = mOutConfigW[19:16]; 
assign MEMC4_data_out_ctx2 = mDataFromMem[159:128]; 
assign mDataToMem[159:128] = MEMC4_data_in_ctx1; 
assign globalDataOut[159:128] = MEMC4_data_to_Core; 
assign MEMC4_valid_ctx1 = valid1[4:4]; 
assign MEMC4_write_en_ctx1 = WEn1[4:4]; 
assign MEMC4_stride_ctx1 = stride1[4:4]; 
assign MEMC4_start_addr_ctx1 = startAddr1[29:24]; 
assign MEMC4_burst_count_ctx1 = count1[34:28]; 
assign mAddr1[29:24] = MEMC4_addr_out_ctx1; 
assign mEn1[4:4] = MEMC4_mem_en_ctx1; 
assign mWEn1[4:4] = MEMC4_write_mem_en_ctx1; 
assign MEMC4_valid_ctx2 = valid2[4:4]; 
assign MEMC4_write_en_ctx2 = WEn2[4:4]; 
assign MEMC4_stride_ctx2 = stride2[4:4]; 
assign MEMC4_start_addr_ctx2 = startAddr2[29:24]; 
assign mAddr2[29:24] = MEMC4_addr_out_ctx2; 
assign MEMC4_burst_count_ctx2 = count2[34:28]; 
assign mEn2[4:4] = MEMC4_mem_en_ctx2; 
assign mWEn2[4:4] = MEMC4_write_mem_en_ctx2; 
wire [31:0] MEMOCMux5_inw1;
wire [31:0] MEMOCMux5_inw2;
wire [31:0] MEMOCMux5_inw3;
wire [31:0] MEMOCMux5_inw4;
wire [31:0] MEMOCMux5_inw5;
wire [31:0] MEMOCMux5_inw6;
wire [31:0] MEMOCMux5_inw7;
wire [31:0] MEMOCMux5_inw8;
wire [31:0] MEMOCMux5_inw9;
wire [31:0] MEMOCMux5_inw10;
wire [31:0] MEMOCMux5_outw1;
wire [3:0] MEMOCMux5_selw;
HA_10IM MEMOCMux5 (
.DataIn_1(MEMOCMux5_inw1),
.DataIn_2(MEMOCMux5_inw2),
.DataIn_3(MEMOCMux5_inw3),
.DataIn_4(MEMOCMux5_inw4),
.DataIn_5(MEMOCMux5_inw5),
.DataIn_6(MEMOCMux5_inw6),
.DataIn_7(MEMOCMux5_inw7),
.DataIn_8(MEMOCMux5_inw8),
.DataIn_9(MEMOCMux5_inw9),
.DataIn_10(MEMOCMux5_inw10),
.DataOut_1(MEMOCMux5_outw1),
.sel(MEMOCMux5_selw));
defparam MEMOCMux5.Mux_BW = 32;
assign MEMC5_data_from_Core = MEMOCMux5_outw1;
assign MEMOCMux5_inw1 = dataOutW[31:0]; 
assign MEMOCMux5_inw2 = dataOutW[63:32]; 
assign MEMOCMux5_inw3 = dataOutW[95:64]; 
assign MEMOCMux5_inw4 = dataOutW[127:96]; 
assign MEMOCMux5_inw5 = dataOutW[159:128]; 
assign MEMOCMux5_inw6 = dataOutW[191:160]; 
assign MEMOCMux5_inw7 = dataOutW[223:192]; 
assign MEMOCMux5_inw8 = dataOutW[255:224]; 
assign MEMOCMux5_inw9 = dataOutW[287:256]; 
assign MEMOCMux5_inw10 = globalDataIn[191:160]; 
assign MEMOCMux5_selw = mOutConfigW[23:20]; 
assign MEMC5_data_out_ctx2 = mDataFromMem[191:160]; 
assign mDataToMem[191:160] = MEMC5_data_in_ctx1; 
assign globalDataOut[191:160] = MEMC5_data_to_Core; 
assign MEMC5_valid_ctx1 = valid1[5:5]; 
assign MEMC5_write_en_ctx1 = WEn1[5:5]; 
assign MEMC5_stride_ctx1 = stride1[5:5]; 
assign MEMC5_start_addr_ctx1 = startAddr1[35:30]; 
assign MEMC5_burst_count_ctx1 = count1[41:35]; 
assign mAddr1[35:30] = MEMC5_addr_out_ctx1; 
assign mEn1[5:5] = MEMC5_mem_en_ctx1; 
assign mWEn1[5:5] = MEMC5_write_mem_en_ctx1; 
assign MEMC5_valid_ctx2 = valid2[5:5]; 
assign MEMC5_write_en_ctx2 = WEn2[5:5]; 
assign MEMC5_stride_ctx2 = stride2[5:5]; 
assign MEMC5_start_addr_ctx2 = startAddr2[35:30]; 
assign mAddr2[35:30] = MEMC5_addr_out_ctx2; 
assign MEMC5_burst_count_ctx2 = count2[41:35]; 
assign mEn2[5:5] = MEMC5_mem_en_ctx2; 
assign mWEn2[5:5] = MEMC5_write_mem_en_ctx2; 
wire [31:0] MEMOCMux6_inw1;
wire [31:0] MEMOCMux6_inw2;
wire [31:0] MEMOCMux6_inw3;
wire [31:0] MEMOCMux6_inw4;
wire [31:0] MEMOCMux6_inw5;
wire [31:0] MEMOCMux6_inw6;
wire [31:0] MEMOCMux6_inw7;
wire [31:0] MEMOCMux6_inw8;
wire [31:0] MEMOCMux6_inw9;
wire [31:0] MEMOCMux6_inw10;
wire [31:0] MEMOCMux6_outw1;
wire [3:0] MEMOCMux6_selw;
HA_10IM MEMOCMux6 (
.DataIn_1(MEMOCMux6_inw1),
.DataIn_2(MEMOCMux6_inw2),
.DataIn_3(MEMOCMux6_inw3),
.DataIn_4(MEMOCMux6_inw4),
.DataIn_5(MEMOCMux6_inw5),
.DataIn_6(MEMOCMux6_inw6),
.DataIn_7(MEMOCMux6_inw7),
.DataIn_8(MEMOCMux6_inw8),
.DataIn_9(MEMOCMux6_inw9),
.DataIn_10(MEMOCMux6_inw10),
.DataOut_1(MEMOCMux6_outw1),
.sel(MEMOCMux6_selw));
defparam MEMOCMux6.Mux_BW = 32;
assign MEMC6_data_from_Core = MEMOCMux6_outw1;
assign MEMOCMux6_inw1 = dataOutW[31:0]; 
assign MEMOCMux6_inw2 = dataOutW[63:32]; 
assign MEMOCMux6_inw3 = dataOutW[95:64]; 
assign MEMOCMux6_inw4 = dataOutW[127:96]; 
assign MEMOCMux6_inw5 = dataOutW[159:128]; 
assign MEMOCMux6_inw6 = dataOutW[191:160]; 
assign MEMOCMux6_inw7 = dataOutW[223:192]; 
assign MEMOCMux6_inw8 = dataOutW[255:224]; 
assign MEMOCMux6_inw9 = dataOutW[287:256]; 
assign MEMOCMux6_inw10 = globalDataIn[223:192]; 
assign MEMOCMux6_selw = mOutConfigW[27:24]; 
assign MEMC6_data_out_ctx2 = mDataFromMem[223:192]; 
assign mDataToMem[223:192] = MEMC6_data_in_ctx1; 
assign globalDataOut[223:192] = MEMC6_data_to_Core; 
assign MEMC6_valid_ctx1 = valid1[6:6]; 
assign MEMC6_write_en_ctx1 = WEn1[6:6]; 
assign MEMC6_stride_ctx1 = stride1[6:6]; 
assign MEMC6_start_addr_ctx1 = startAddr1[41:36]; 
assign MEMC6_burst_count_ctx1 = count1[48:42]; 
assign mAddr1[41:36] = MEMC6_addr_out_ctx1; 
assign mEn1[6:6] = MEMC6_mem_en_ctx1; 
assign mWEn1[6:6] = MEMC6_write_mem_en_ctx1; 
assign MEMC6_valid_ctx2 = valid2[6:6]; 
assign MEMC6_write_en_ctx2 = WEn2[6:6]; 
assign MEMC6_stride_ctx2 = stride2[6:6]; 
assign MEMC6_start_addr_ctx2 = startAddr2[41:36]; 
assign mAddr2[41:36] = MEMC6_addr_out_ctx2; 
assign MEMC6_burst_count_ctx2 = count2[48:42]; 
assign mEn2[6:6] = MEMC6_mem_en_ctx2; 
assign mWEn2[6:6] = MEMC6_write_mem_en_ctx2; 
wire [31:0] MEMOCMux7_inw1;
wire [31:0] MEMOCMux7_inw2;
wire [31:0] MEMOCMux7_inw3;
wire [31:0] MEMOCMux7_inw4;
wire [31:0] MEMOCMux7_inw5;
wire [31:0] MEMOCMux7_inw6;
wire [31:0] MEMOCMux7_inw7;
wire [31:0] MEMOCMux7_inw8;
wire [31:0] MEMOCMux7_inw9;
wire [31:0] MEMOCMux7_inw10;
wire [31:0] MEMOCMux7_outw1;
wire [3:0] MEMOCMux7_selw;
HA_10IM MEMOCMux7 (
.DataIn_1(MEMOCMux7_inw1),
.DataIn_2(MEMOCMux7_inw2),
.DataIn_3(MEMOCMux7_inw3),
.DataIn_4(MEMOCMux7_inw4),
.DataIn_5(MEMOCMux7_inw5),
.DataIn_6(MEMOCMux7_inw6),
.DataIn_7(MEMOCMux7_inw7),
.DataIn_8(MEMOCMux7_inw8),
.DataIn_9(MEMOCMux7_inw9),
.DataIn_10(MEMOCMux7_inw10),
.DataOut_1(MEMOCMux7_outw1),
.sel(MEMOCMux7_selw));
defparam MEMOCMux7.Mux_BW = 32;
assign MEMC7_data_from_Core = MEMOCMux7_outw1;
assign MEMOCMux7_inw1 = dataOutW[31:0]; 
assign MEMOCMux7_inw2 = dataOutW[63:32]; 
assign MEMOCMux7_inw3 = dataOutW[95:64]; 
assign MEMOCMux7_inw4 = dataOutW[127:96]; 
assign MEMOCMux7_inw5 = dataOutW[159:128]; 
assign MEMOCMux7_inw6 = dataOutW[191:160]; 
assign MEMOCMux7_inw7 = dataOutW[223:192]; 
assign MEMOCMux7_inw8 = dataOutW[255:224]; 
assign MEMOCMux7_inw9 = dataOutW[287:256]; 
assign MEMOCMux7_inw10 = globalDataIn[255:224]; 
assign MEMOCMux7_selw = mOutConfigW[31:28]; 
assign MEMC7_data_out_ctx2 = mDataFromMem[255:224]; 
assign mDataToMem[255:224] = MEMC7_data_in_ctx1; 
assign globalDataOut[255:224] = MEMC7_data_to_Core; 
assign MEMC7_valid_ctx1 = valid1[7:7]; 
assign MEMC7_write_en_ctx1 = WEn1[7:7]; 
assign MEMC7_stride_ctx1 = stride1[7:7]; 
assign MEMC7_start_addr_ctx1 = startAddr1[47:42]; 
assign MEMC7_burst_count_ctx1 = count1[55:49]; 
assign mAddr1[47:42] = MEMC7_addr_out_ctx1; 
assign mEn1[7:7] = MEMC7_mem_en_ctx1; 
assign mWEn1[7:7] = MEMC7_write_mem_en_ctx1; 
assign MEMC7_valid_ctx2 = valid2[7:7]; 
assign MEMC7_write_en_ctx2 = WEn2[7:7]; 
assign MEMC7_stride_ctx2 = stride2[7:7]; 
assign MEMC7_start_addr_ctx2 = startAddr2[47:42]; 
assign mAddr2[47:42] = MEMC7_addr_out_ctx2; 
assign MEMC7_burst_count_ctx2 = count2[55:49]; 
assign mEn2[7:7] = MEMC7_mem_en_ctx2; 
assign mWEn2[7:7] = MEMC7_write_mem_en_ctx2; 
wire [31:0] MEMOCMux8_inw1;
wire [31:0] MEMOCMux8_inw2;
wire [31:0] MEMOCMux8_inw3;
wire [31:0] MEMOCMux8_inw4;
wire [31:0] MEMOCMux8_inw5;
wire [31:0] MEMOCMux8_inw6;
wire [31:0] MEMOCMux8_inw7;
wire [31:0] MEMOCMux8_inw8;
wire [31:0] MEMOCMux8_inw9;
wire [31:0] MEMOCMux8_inw10;
wire [31:0] MEMOCMux8_outw1;
wire [3:0] MEMOCMux8_selw;
HA_10IM MEMOCMux8 (
.DataIn_1(MEMOCMux8_inw1),
.DataIn_2(MEMOCMux8_inw2),
.DataIn_3(MEMOCMux8_inw3),
.DataIn_4(MEMOCMux8_inw4),
.DataIn_5(MEMOCMux8_inw5),
.DataIn_6(MEMOCMux8_inw6),
.DataIn_7(MEMOCMux8_inw7),
.DataIn_8(MEMOCMux8_inw8),
.DataIn_9(MEMOCMux8_inw9),
.DataIn_10(MEMOCMux8_inw10),
.DataOut_1(MEMOCMux8_outw1),
.sel(MEMOCMux8_selw));
defparam MEMOCMux8.Mux_BW = 32;
assign MEMC8_data_from_Core = MEMOCMux8_outw1;
assign MEMOCMux8_inw1 = dataOutW[31:0]; 
assign MEMOCMux8_inw2 = dataOutW[63:32]; 
assign MEMOCMux8_inw3 = dataOutW[95:64]; 
assign MEMOCMux8_inw4 = dataOutW[127:96]; 
assign MEMOCMux8_inw5 = dataOutW[159:128]; 
assign MEMOCMux8_inw6 = dataOutW[191:160]; 
assign MEMOCMux8_inw7 = dataOutW[223:192]; 
assign MEMOCMux8_inw8 = dataOutW[255:224]; 
assign MEMOCMux8_inw9 = dataOutW[287:256]; 
assign MEMOCMux8_inw10 = globalDataIn[287:256]; 
assign MEMOCMux8_selw = mOutConfigW[35:32]; 
assign MEMC8_data_out_ctx2 = mDataFromMem[287:256]; 
assign mDataToMem[287:256] = MEMC8_data_in_ctx1; 
assign globalDataOut[287:256] = MEMC8_data_to_Core; 
assign MEMC8_valid_ctx1 = valid1[8:8]; 
assign MEMC8_write_en_ctx1 = WEn1[8:8]; 
assign MEMC8_stride_ctx1 = stride1[8:8]; 
assign MEMC8_start_addr_ctx1 = startAddr1[53:48]; 
assign MEMC8_burst_count_ctx1 = count1[62:56]; 
assign mAddr1[53:48] = MEMC8_addr_out_ctx1; 
assign mEn1[8:8] = MEMC8_mem_en_ctx1; 
assign mWEn1[8:8] = MEMC8_write_mem_en_ctx1; 
assign MEMC8_valid_ctx2 = valid2[8:8]; 
assign MEMC8_write_en_ctx2 = WEn2[8:8]; 
assign MEMC8_stride_ctx2 = stride2[8:8]; 
assign MEMC8_start_addr_ctx2 = startAddr2[53:48]; 
assign mAddr2[53:48] = MEMC8_addr_out_ctx2; 
assign MEMC8_burst_count_ctx2 = count2[62:56]; 
assign mEn2[8:8] = MEMC8_mem_en_ctx2; 
assign mWEn2[8:8] = MEMC8_write_mem_en_ctx2; 
wire [31:0] MEMOCMux9_inw1;
wire [31:0] MEMOCMux9_inw2;
wire [31:0] MEMOCMux9_inw3;
wire [31:0] MEMOCMux9_inw4;
wire [31:0] MEMOCMux9_inw5;
wire [31:0] MEMOCMux9_inw6;
wire [31:0] MEMOCMux9_inw7;
wire [31:0] MEMOCMux9_inw8;
wire [31:0] MEMOCMux9_inw9;
wire [31:0] MEMOCMux9_inw10;
wire [31:0] MEMOCMux9_outw1;
wire [3:0] MEMOCMux9_selw;
HA_10IM MEMOCMux9 (
.DataIn_1(MEMOCMux9_inw1),
.DataIn_2(MEMOCMux9_inw2),
.DataIn_3(MEMOCMux9_inw3),
.DataIn_4(MEMOCMux9_inw4),
.DataIn_5(MEMOCMux9_inw5),
.DataIn_6(MEMOCMux9_inw6),
.DataIn_7(MEMOCMux9_inw7),
.DataIn_8(MEMOCMux9_inw8),
.DataIn_9(MEMOCMux9_inw9),
.DataIn_10(MEMOCMux9_inw10),
.DataOut_1(MEMOCMux9_outw1),
.sel(MEMOCMux9_selw));
defparam MEMOCMux9.Mux_BW = 32;
assign MEMC9_data_from_Core = MEMOCMux9_outw1;
assign MEMOCMux9_inw1 = dataOutW[31:0]; 
assign MEMOCMux9_inw2 = dataOutW[63:32]; 
assign MEMOCMux9_inw3 = dataOutW[95:64]; 
assign MEMOCMux9_inw4 = dataOutW[127:96]; 
assign MEMOCMux9_inw5 = dataOutW[159:128]; 
assign MEMOCMux9_inw6 = dataOutW[191:160]; 
assign MEMOCMux9_inw7 = dataOutW[223:192]; 
assign MEMOCMux9_inw8 = dataOutW[255:224]; 
assign MEMOCMux9_inw9 = dataOutW[287:256]; 
assign MEMOCMux9_inw10 = globalDataIn[319:288]; 
assign MEMOCMux9_selw = mOutConfigW[39:36]; 
assign MEMC9_data_out_ctx2 = mDataFromMem[319:288]; 
assign mDataToMem[319:288] = MEMC9_data_in_ctx1; 
assign globalDataOut[319:288] = MEMC9_data_to_Core; 
assign MEMC9_valid_ctx1 = valid1[9:9]; 
assign MEMC9_write_en_ctx1 = WEn1[9:9]; 
assign MEMC9_stride_ctx1 = stride1[9:9]; 
assign MEMC9_start_addr_ctx1 = startAddr1[59:54]; 
assign MEMC9_burst_count_ctx1 = count1[69:63]; 
assign mAddr1[59:54] = MEMC9_addr_out_ctx1; 
assign mEn1[9:9] = MEMC9_mem_en_ctx1; 
assign mWEn1[9:9] = MEMC9_write_mem_en_ctx1; 
assign MEMC9_valid_ctx2 = valid2[9:9]; 
assign MEMC9_write_en_ctx2 = WEn2[9:9]; 
assign MEMC9_stride_ctx2 = stride2[9:9]; 
assign MEMC9_start_addr_ctx2 = startAddr2[59:54]; 
assign mAddr2[59:54] = MEMC9_addr_out_ctx2; 
assign MEMC9_burst_count_ctx2 = count2[69:63]; 
assign mEn2[9:9] = MEMC9_mem_en_ctx2; 
assign mWEn2[9:9] = MEMC9_write_mem_en_ctx2; 
wire [31:0] MEMOCMux10_inw1;
wire [31:0] MEMOCMux10_inw2;
wire [31:0] MEMOCMux10_inw3;
wire [31:0] MEMOCMux10_inw4;
wire [31:0] MEMOCMux10_inw5;
wire [31:0] MEMOCMux10_inw6;
wire [31:0] MEMOCMux10_inw7;
wire [31:0] MEMOCMux10_inw8;
wire [31:0] MEMOCMux10_inw9;
wire [31:0] MEMOCMux10_inw10;
wire [31:0] MEMOCMux10_outw1;
wire [3:0] MEMOCMux10_selw;
HA_10IM MEMOCMux10 (
.DataIn_1(MEMOCMux10_inw1),
.DataIn_2(MEMOCMux10_inw2),
.DataIn_3(MEMOCMux10_inw3),
.DataIn_4(MEMOCMux10_inw4),
.DataIn_5(MEMOCMux10_inw5),
.DataIn_6(MEMOCMux10_inw6),
.DataIn_7(MEMOCMux10_inw7),
.DataIn_8(MEMOCMux10_inw8),
.DataIn_9(MEMOCMux10_inw9),
.DataIn_10(MEMOCMux10_inw10),
.DataOut_1(MEMOCMux10_outw1),
.sel(MEMOCMux10_selw));
defparam MEMOCMux10.Mux_BW = 32;
assign MEMC10_data_from_Core = MEMOCMux10_outw1;
assign MEMOCMux10_inw1 = dataOutW[31:0]; 
assign MEMOCMux10_inw2 = dataOutW[63:32]; 
assign MEMOCMux10_inw3 = dataOutW[95:64]; 
assign MEMOCMux10_inw4 = dataOutW[127:96]; 
assign MEMOCMux10_inw5 = dataOutW[159:128]; 
assign MEMOCMux10_inw6 = dataOutW[191:160]; 
assign MEMOCMux10_inw7 = dataOutW[223:192]; 
assign MEMOCMux10_inw8 = dataOutW[255:224]; 
assign MEMOCMux10_inw9 = dataOutW[287:256]; 
assign MEMOCMux10_inw10 = globalDataIn[351:320]; 
assign MEMOCMux10_selw = mOutConfigW[43:40]; 
assign MEMC10_data_out_ctx2 = mDataFromMem[351:320]; 
assign mDataToMem[351:320] = MEMC10_data_in_ctx1; 
assign globalDataOut[351:320] = MEMC10_data_to_Core; 
assign MEMC10_valid_ctx1 = valid1[10:10]; 
assign MEMC10_write_en_ctx1 = WEn1[10:10]; 
assign MEMC10_stride_ctx1 = stride1[10:10]; 
assign MEMC10_start_addr_ctx1 = startAddr1[65:60]; 
assign MEMC10_burst_count_ctx1 = count1[76:70]; 
assign mAddr1[65:60] = MEMC10_addr_out_ctx1; 
assign mEn1[10:10] = MEMC10_mem_en_ctx1; 
assign mWEn1[10:10] = MEMC10_write_mem_en_ctx1; 
assign MEMC10_valid_ctx2 = valid2[10:10]; 
assign MEMC10_write_en_ctx2 = WEn2[10:10]; 
assign MEMC10_stride_ctx2 = stride2[10:10]; 
assign MEMC10_start_addr_ctx2 = startAddr2[65:60]; 
assign mAddr2[65:60] = MEMC10_addr_out_ctx2; 
assign MEMC10_burst_count_ctx2 = count2[76:70]; 
assign mEn2[10:10] = MEMC10_mem_en_ctx2; 
assign mWEn2[10:10] = MEMC10_write_mem_en_ctx2; 
wire [31:0] MEMOCMux11_inw1;
wire [31:0] MEMOCMux11_inw2;
wire [31:0] MEMOCMux11_inw3;
wire [31:0] MEMOCMux11_inw4;
wire [31:0] MEMOCMux11_inw5;
wire [31:0] MEMOCMux11_inw6;
wire [31:0] MEMOCMux11_inw7;
wire [31:0] MEMOCMux11_inw8;
wire [31:0] MEMOCMux11_inw9;
wire [31:0] MEMOCMux11_inw10;
wire [31:0] MEMOCMux11_outw1;
wire [3:0] MEMOCMux11_selw;
HA_10IM MEMOCMux11 (
.DataIn_1(MEMOCMux11_inw1),
.DataIn_2(MEMOCMux11_inw2),
.DataIn_3(MEMOCMux11_inw3),
.DataIn_4(MEMOCMux11_inw4),
.DataIn_5(MEMOCMux11_inw5),
.DataIn_6(MEMOCMux11_inw6),
.DataIn_7(MEMOCMux11_inw7),
.DataIn_8(MEMOCMux11_inw8),
.DataIn_9(MEMOCMux11_inw9),
.DataIn_10(MEMOCMux11_inw10),
.DataOut_1(MEMOCMux11_outw1),
.sel(MEMOCMux11_selw));
defparam MEMOCMux11.Mux_BW = 32;
assign MEMC11_data_from_Core = MEMOCMux11_outw1;
assign MEMOCMux11_inw1 = dataOutW[31:0]; 
assign MEMOCMux11_inw2 = dataOutW[63:32]; 
assign MEMOCMux11_inw3 = dataOutW[95:64]; 
assign MEMOCMux11_inw4 = dataOutW[127:96]; 
assign MEMOCMux11_inw5 = dataOutW[159:128]; 
assign MEMOCMux11_inw6 = dataOutW[191:160]; 
assign MEMOCMux11_inw7 = dataOutW[223:192]; 
assign MEMOCMux11_inw8 = dataOutW[255:224]; 
assign MEMOCMux11_inw9 = dataOutW[287:256]; 
assign MEMOCMux11_inw10 = globalDataIn[383:352]; 
assign MEMOCMux11_selw = mOutConfigW[47:44]; 
assign MEMC11_data_out_ctx2 = mDataFromMem[383:352]; 
assign mDataToMem[383:352] = MEMC11_data_in_ctx1; 
assign globalDataOut[383:352] = MEMC11_data_to_Core; 
assign MEMC11_valid_ctx1 = valid1[11:11]; 
assign MEMC11_write_en_ctx1 = WEn1[11:11]; 
assign MEMC11_stride_ctx1 = stride1[11:11]; 
assign MEMC11_start_addr_ctx1 = startAddr1[71:66]; 
assign MEMC11_burst_count_ctx1 = count1[83:77]; 
assign mAddr1[71:66] = MEMC11_addr_out_ctx1; 
assign mEn1[11:11] = MEMC11_mem_en_ctx1; 
assign mWEn1[11:11] = MEMC11_write_mem_en_ctx1; 
assign MEMC11_valid_ctx2 = valid2[11:11]; 
assign MEMC11_write_en_ctx2 = WEn2[11:11]; 
assign MEMC11_stride_ctx2 = stride2[11:11]; 
assign MEMC11_start_addr_ctx2 = startAddr2[71:66]; 
assign mAddr2[71:66] = MEMC11_addr_out_ctx2; 
assign MEMC11_burst_count_ctx2 = count2[83:77]; 
assign mEn2[11:11] = MEMC11_mem_en_ctx2; 
assign mWEn2[11:11] = MEMC11_write_mem_en_ctx2; 
wire [31:0] MEMOCMux12_inw1;
wire [31:0] MEMOCMux12_inw2;
wire [31:0] MEMOCMux12_inw3;
wire [31:0] MEMOCMux12_inw4;
wire [31:0] MEMOCMux12_inw5;
wire [31:0] MEMOCMux12_inw6;
wire [31:0] MEMOCMux12_inw7;
wire [31:0] MEMOCMux12_inw8;
wire [31:0] MEMOCMux12_inw9;
wire [31:0] MEMOCMux12_inw10;
wire [31:0] MEMOCMux12_outw1;
wire [3:0] MEMOCMux12_selw;
HA_10IM MEMOCMux12 (
.DataIn_1(MEMOCMux12_inw1),
.DataIn_2(MEMOCMux12_inw2),
.DataIn_3(MEMOCMux12_inw3),
.DataIn_4(MEMOCMux12_inw4),
.DataIn_5(MEMOCMux12_inw5),
.DataIn_6(MEMOCMux12_inw6),
.DataIn_7(MEMOCMux12_inw7),
.DataIn_8(MEMOCMux12_inw8),
.DataIn_9(MEMOCMux12_inw9),
.DataIn_10(MEMOCMux12_inw10),
.DataOut_1(MEMOCMux12_outw1),
.sel(MEMOCMux12_selw));
defparam MEMOCMux12.Mux_BW = 32;
assign MEMC12_data_from_Core = MEMOCMux12_outw1;
assign MEMOCMux12_inw1 = dataOutW[31:0]; 
assign MEMOCMux12_inw2 = dataOutW[63:32]; 
assign MEMOCMux12_inw3 = dataOutW[95:64]; 
assign MEMOCMux12_inw4 = dataOutW[127:96]; 
assign MEMOCMux12_inw5 = dataOutW[159:128]; 
assign MEMOCMux12_inw6 = dataOutW[191:160]; 
assign MEMOCMux12_inw7 = dataOutW[223:192]; 
assign MEMOCMux12_inw8 = dataOutW[255:224]; 
assign MEMOCMux12_inw9 = dataOutW[287:256]; 
assign MEMOCMux12_inw10 = globalDataIn[415:384]; 
assign MEMOCMux12_selw = mOutConfigW[51:48]; 
assign MEMC12_data_out_ctx2 = mDataFromMem[415:384]; 
assign mDataToMem[415:384] = MEMC12_data_in_ctx1; 
assign globalDataOut[415:384] = MEMC12_data_to_Core; 
assign MEMC12_valid_ctx1 = valid1[12:12]; 
assign MEMC12_write_en_ctx1 = WEn1[12:12]; 
assign MEMC12_stride_ctx1 = stride1[12:12]; 
assign MEMC12_start_addr_ctx1 = startAddr1[77:72]; 
assign MEMC12_burst_count_ctx1 = count1[90:84]; 
assign mAddr1[77:72] = MEMC12_addr_out_ctx1; 
assign mEn1[12:12] = MEMC12_mem_en_ctx1; 
assign mWEn1[12:12] = MEMC12_write_mem_en_ctx1; 
assign MEMC12_valid_ctx2 = valid2[12:12]; 
assign MEMC12_write_en_ctx2 = WEn2[12:12]; 
assign MEMC12_stride_ctx2 = stride2[12:12]; 
assign MEMC12_start_addr_ctx2 = startAddr2[77:72]; 
assign mAddr2[77:72] = MEMC12_addr_out_ctx2; 
assign MEMC12_burst_count_ctx2 = count2[90:84]; 
assign mEn2[12:12] = MEMC12_mem_en_ctx2; 
assign mWEn2[12:12] = MEMC12_write_mem_en_ctx2; 
wire [31:0] MEMOCMux13_inw1;
wire [31:0] MEMOCMux13_inw2;
wire [31:0] MEMOCMux13_inw3;
wire [31:0] MEMOCMux13_inw4;
wire [31:0] MEMOCMux13_inw5;
wire [31:0] MEMOCMux13_inw6;
wire [31:0] MEMOCMux13_inw7;
wire [31:0] MEMOCMux13_inw8;
wire [31:0] MEMOCMux13_inw9;
wire [31:0] MEMOCMux13_inw10;
wire [31:0] MEMOCMux13_outw1;
wire [3:0] MEMOCMux13_selw;
HA_10IM MEMOCMux13 (
.DataIn_1(MEMOCMux13_inw1),
.DataIn_2(MEMOCMux13_inw2),
.DataIn_3(MEMOCMux13_inw3),
.DataIn_4(MEMOCMux13_inw4),
.DataIn_5(MEMOCMux13_inw5),
.DataIn_6(MEMOCMux13_inw6),
.DataIn_7(MEMOCMux13_inw7),
.DataIn_8(MEMOCMux13_inw8),
.DataIn_9(MEMOCMux13_inw9),
.DataIn_10(MEMOCMux13_inw10),
.DataOut_1(MEMOCMux13_outw1),
.sel(MEMOCMux13_selw));
defparam MEMOCMux13.Mux_BW = 32;
assign MEMC13_data_from_Core = MEMOCMux13_outw1;
assign MEMOCMux13_inw1 = dataOutW[31:0]; 
assign MEMOCMux13_inw2 = dataOutW[63:32]; 
assign MEMOCMux13_inw3 = dataOutW[95:64]; 
assign MEMOCMux13_inw4 = dataOutW[127:96]; 
assign MEMOCMux13_inw5 = dataOutW[159:128]; 
assign MEMOCMux13_inw6 = dataOutW[191:160]; 
assign MEMOCMux13_inw7 = dataOutW[223:192]; 
assign MEMOCMux13_inw8 = dataOutW[255:224]; 
assign MEMOCMux13_inw9 = dataOutW[287:256]; 
assign MEMOCMux13_inw10 = globalDataIn[447:416]; 
assign MEMOCMux13_selw = mOutConfigW[55:52]; 
assign MEMC13_data_out_ctx2 = mDataFromMem[447:416]; 
assign mDataToMem[447:416] = MEMC13_data_in_ctx1; 
assign globalDataOut[447:416] = MEMC13_data_to_Core; 
assign MEMC13_valid_ctx1 = valid1[13:13]; 
assign MEMC13_write_en_ctx1 = WEn1[13:13]; 
assign MEMC13_stride_ctx1 = stride1[13:13]; 
assign MEMC13_start_addr_ctx1 = startAddr1[83:78]; 
assign MEMC13_burst_count_ctx1 = count1[97:91]; 
assign mAddr1[83:78] = MEMC13_addr_out_ctx1; 
assign mEn1[13:13] = MEMC13_mem_en_ctx1; 
assign mWEn1[13:13] = MEMC13_write_mem_en_ctx1; 
assign MEMC13_valid_ctx2 = valid2[13:13]; 
assign MEMC13_write_en_ctx2 = WEn2[13:13]; 
assign MEMC13_stride_ctx2 = stride2[13:13]; 
assign MEMC13_start_addr_ctx2 = startAddr2[83:78]; 
assign mAddr2[83:78] = MEMC13_addr_out_ctx2; 
assign MEMC13_burst_count_ctx2 = count2[97:91]; 
assign mEn2[13:13] = MEMC13_mem_en_ctx2; 
assign mWEn2[13:13] = MEMC13_write_mem_en_ctx2; 
wire [31:0] MEMOCMux14_inw1;
wire [31:0] MEMOCMux14_inw2;
wire [31:0] MEMOCMux14_inw3;
wire [31:0] MEMOCMux14_inw4;
wire [31:0] MEMOCMux14_inw5;
wire [31:0] MEMOCMux14_inw6;
wire [31:0] MEMOCMux14_inw7;
wire [31:0] MEMOCMux14_inw8;
wire [31:0] MEMOCMux14_inw9;
wire [31:0] MEMOCMux14_inw10;
wire [31:0] MEMOCMux14_outw1;
wire [3:0] MEMOCMux14_selw;
HA_10IM MEMOCMux14 (
.DataIn_1(MEMOCMux14_inw1),
.DataIn_2(MEMOCMux14_inw2),
.DataIn_3(MEMOCMux14_inw3),
.DataIn_4(MEMOCMux14_inw4),
.DataIn_5(MEMOCMux14_inw5),
.DataIn_6(MEMOCMux14_inw6),
.DataIn_7(MEMOCMux14_inw7),
.DataIn_8(MEMOCMux14_inw8),
.DataIn_9(MEMOCMux14_inw9),
.DataIn_10(MEMOCMux14_inw10),
.DataOut_1(MEMOCMux14_outw1),
.sel(MEMOCMux14_selw));
defparam MEMOCMux14.Mux_BW = 32;
assign MEMC14_data_from_Core = MEMOCMux14_outw1;
assign MEMOCMux14_inw1 = dataOutW[31:0]; 
assign MEMOCMux14_inw2 = dataOutW[63:32]; 
assign MEMOCMux14_inw3 = dataOutW[95:64]; 
assign MEMOCMux14_inw4 = dataOutW[127:96]; 
assign MEMOCMux14_inw5 = dataOutW[159:128]; 
assign MEMOCMux14_inw6 = dataOutW[191:160]; 
assign MEMOCMux14_inw7 = dataOutW[223:192]; 
assign MEMOCMux14_inw8 = dataOutW[255:224]; 
assign MEMOCMux14_inw9 = dataOutW[287:256]; 
assign MEMOCMux14_inw10 = globalDataIn[479:448]; 
assign MEMOCMux14_selw = mOutConfigW[59:56]; 
assign MEMC14_data_out_ctx2 = mDataFromMem[479:448]; 
assign mDataToMem[479:448] = MEMC14_data_in_ctx1; 
assign globalDataOut[479:448] = MEMC14_data_to_Core; 
assign MEMC14_valid_ctx1 = valid1[14:14]; 
assign MEMC14_write_en_ctx1 = WEn1[14:14]; 
assign MEMC14_stride_ctx1 = stride1[14:14]; 
assign MEMC14_start_addr_ctx1 = startAddr1[89:84]; 
assign MEMC14_burst_count_ctx1 = count1[104:98]; 
assign mAddr1[89:84] = MEMC14_addr_out_ctx1; 
assign mEn1[14:14] = MEMC14_mem_en_ctx1; 
assign mWEn1[14:14] = MEMC14_write_mem_en_ctx1; 
assign MEMC14_valid_ctx2 = valid2[14:14]; 
assign MEMC14_write_en_ctx2 = WEn2[14:14]; 
assign MEMC14_stride_ctx2 = stride2[14:14]; 
assign MEMC14_start_addr_ctx2 = startAddr2[89:84]; 
assign mAddr2[89:84] = MEMC14_addr_out_ctx2; 
assign MEMC14_burst_count_ctx2 = count2[104:98]; 
assign mEn2[14:14] = MEMC14_mem_en_ctx2; 
assign mWEn2[14:14] = MEMC14_write_mem_en_ctx2; 
wire [31:0] MEMOCMux15_inw1;
wire [31:0] MEMOCMux15_inw2;
wire [31:0] MEMOCMux15_inw3;
wire [31:0] MEMOCMux15_inw4;
wire [31:0] MEMOCMux15_inw5;
wire [31:0] MEMOCMux15_inw6;
wire [31:0] MEMOCMux15_inw7;
wire [31:0] MEMOCMux15_inw8;
wire [31:0] MEMOCMux15_inw9;
wire [31:0] MEMOCMux15_inw10;
wire [31:0] MEMOCMux15_outw1;
wire [3:0] MEMOCMux15_selw;
HA_10IM MEMOCMux15 (
.DataIn_1(MEMOCMux15_inw1),
.DataIn_2(MEMOCMux15_inw2),
.DataIn_3(MEMOCMux15_inw3),
.DataIn_4(MEMOCMux15_inw4),
.DataIn_5(MEMOCMux15_inw5),
.DataIn_6(MEMOCMux15_inw6),
.DataIn_7(MEMOCMux15_inw7),
.DataIn_8(MEMOCMux15_inw8),
.DataIn_9(MEMOCMux15_inw9),
.DataIn_10(MEMOCMux15_inw10),
.DataOut_1(MEMOCMux15_outw1),
.sel(MEMOCMux15_selw));
defparam MEMOCMux15.Mux_BW = 32;
assign MEMC15_data_from_Core = MEMOCMux15_outw1;
assign MEMOCMux15_inw1 = dataOutW[31:0]; 
assign MEMOCMux15_inw2 = dataOutW[63:32]; 
assign MEMOCMux15_inw3 = dataOutW[95:64]; 
assign MEMOCMux15_inw4 = dataOutW[127:96]; 
assign MEMOCMux15_inw5 = dataOutW[159:128]; 
assign MEMOCMux15_inw6 = dataOutW[191:160]; 
assign MEMOCMux15_inw7 = dataOutW[223:192]; 
assign MEMOCMux15_inw8 = dataOutW[255:224]; 
assign MEMOCMux15_inw9 = dataOutW[287:256]; 
assign MEMOCMux15_inw10 = globalDataIn[511:480]; 
assign MEMOCMux15_selw = mOutConfigW[63:60]; 
assign MEMC15_data_out_ctx2 = mDataFromMem[511:480]; 
assign mDataToMem[511:480] = MEMC15_data_in_ctx1; 
assign globalDataOut[511:480] = MEMC15_data_to_Core; 
assign MEMC15_valid_ctx1 = valid1[15:15]; 
assign MEMC15_write_en_ctx1 = WEn1[15:15]; 
assign MEMC15_stride_ctx1 = stride1[15:15]; 
assign MEMC15_start_addr_ctx1 = startAddr1[95:90]; 
assign MEMC15_burst_count_ctx1 = count1[111:105]; 
assign mAddr1[95:90] = MEMC15_addr_out_ctx1; 
assign mEn1[15:15] = MEMC15_mem_en_ctx1; 
assign mWEn1[15:15] = MEMC15_write_mem_en_ctx1; 
assign MEMC15_valid_ctx2 = valid2[15:15]; 
assign MEMC15_write_en_ctx2 = WEn2[15:15]; 
assign MEMC15_stride_ctx2 = stride2[15:15]; 
assign MEMC15_start_addr_ctx2 = startAddr2[95:90]; 
assign mAddr2[95:90] = MEMC15_addr_out_ctx2; 
assign MEMC15_burst_count_ctx2 = count2[111:105]; 
assign mEn2[15:15] = MEMC15_mem_en_ctx2; 
assign mWEn2[15:15] = MEMC15_write_mem_en_ctx2; 
wire [31:0] MEMOCMux16_inw1;
wire [31:0] MEMOCMux16_inw2;
wire [31:0] MEMOCMux16_inw3;
wire [31:0] MEMOCMux16_inw4;
wire [31:0] MEMOCMux16_inw5;
wire [31:0] MEMOCMux16_inw6;
wire [31:0] MEMOCMux16_inw7;
wire [31:0] MEMOCMux16_inw8;
wire [31:0] MEMOCMux16_inw9;
wire [31:0] MEMOCMux16_inw10;
wire [31:0] MEMOCMux16_outw1;
wire [3:0] MEMOCMux16_selw;
HA_10IM MEMOCMux16 (
.DataIn_1(MEMOCMux16_inw1),
.DataIn_2(MEMOCMux16_inw2),
.DataIn_3(MEMOCMux16_inw3),
.DataIn_4(MEMOCMux16_inw4),
.DataIn_5(MEMOCMux16_inw5),
.DataIn_6(MEMOCMux16_inw6),
.DataIn_7(MEMOCMux16_inw7),
.DataIn_8(MEMOCMux16_inw8),
.DataIn_9(MEMOCMux16_inw9),
.DataIn_10(MEMOCMux16_inw10),
.DataOut_1(MEMOCMux16_outw1),
.sel(MEMOCMux16_selw));
defparam MEMOCMux16.Mux_BW = 32;
assign MEMC16_data_from_Core = MEMOCMux16_outw1;
assign MEMOCMux16_inw1 = dataOutW[31:0]; 
assign MEMOCMux16_inw2 = dataOutW[63:32]; 
assign MEMOCMux16_inw3 = dataOutW[95:64]; 
assign MEMOCMux16_inw4 = dataOutW[127:96]; 
assign MEMOCMux16_inw5 = dataOutW[159:128]; 
assign MEMOCMux16_inw6 = dataOutW[191:160]; 
assign MEMOCMux16_inw7 = dataOutW[223:192]; 
assign MEMOCMux16_inw8 = dataOutW[255:224]; 
assign MEMOCMux16_inw9 = dataOutW[287:256]; 
assign MEMOCMux16_inw10 = globalDataIn[543:512]; 
assign MEMOCMux16_selw = mOutConfigW[67:64]; 
assign MEMC16_data_out_ctx2 = mDataFromMem[543:512]; 
assign mDataToMem[543:512] = MEMC16_data_in_ctx1; 
assign globalDataOut[543:512] = MEMC16_data_to_Core; 
assign MEMC16_valid_ctx1 = valid1[16:16]; 
assign MEMC16_write_en_ctx1 = WEn1[16:16]; 
assign MEMC16_stride_ctx1 = stride1[16:16]; 
assign MEMC16_start_addr_ctx1 = startAddr1[101:96]; 
assign MEMC16_burst_count_ctx1 = count1[118:112]; 
assign mAddr1[101:96] = MEMC16_addr_out_ctx1; 
assign mEn1[16:16] = MEMC16_mem_en_ctx1; 
assign mWEn1[16:16] = MEMC16_write_mem_en_ctx1; 
assign MEMC16_valid_ctx2 = valid2[16:16]; 
assign MEMC16_write_en_ctx2 = WEn2[16:16]; 
assign MEMC16_stride_ctx2 = stride2[16:16]; 
assign MEMC16_start_addr_ctx2 = startAddr2[101:96]; 
assign mAddr2[101:96] = MEMC16_addr_out_ctx2; 
assign MEMC16_burst_count_ctx2 = count2[118:112]; 
assign mEn2[16:16] = MEMC16_mem_en_ctx2; 
assign mWEn2[16:16] = MEMC16_write_mem_en_ctx2; 
wire [31:0] MEMOCMux17_inw1;
wire [31:0] MEMOCMux17_inw2;
wire [31:0] MEMOCMux17_inw3;
wire [31:0] MEMOCMux17_inw4;
wire [31:0] MEMOCMux17_inw5;
wire [31:0] MEMOCMux17_inw6;
wire [31:0] MEMOCMux17_inw7;
wire [31:0] MEMOCMux17_inw8;
wire [31:0] MEMOCMux17_inw9;
wire [31:0] MEMOCMux17_inw10;
wire [31:0] MEMOCMux17_outw1;
wire [3:0] MEMOCMux17_selw;
HA_10IM MEMOCMux17 (
.DataIn_1(MEMOCMux17_inw1),
.DataIn_2(MEMOCMux17_inw2),
.DataIn_3(MEMOCMux17_inw3),
.DataIn_4(MEMOCMux17_inw4),
.DataIn_5(MEMOCMux17_inw5),
.DataIn_6(MEMOCMux17_inw6),
.DataIn_7(MEMOCMux17_inw7),
.DataIn_8(MEMOCMux17_inw8),
.DataIn_9(MEMOCMux17_inw9),
.DataIn_10(MEMOCMux17_inw10),
.DataOut_1(MEMOCMux17_outw1),
.sel(MEMOCMux17_selw));
defparam MEMOCMux17.Mux_BW = 32;
assign MEMC17_data_from_Core = MEMOCMux17_outw1;
assign MEMOCMux17_inw1 = dataOutW[31:0]; 
assign MEMOCMux17_inw2 = dataOutW[63:32]; 
assign MEMOCMux17_inw3 = dataOutW[95:64]; 
assign MEMOCMux17_inw4 = dataOutW[127:96]; 
assign MEMOCMux17_inw5 = dataOutW[159:128]; 
assign MEMOCMux17_inw6 = dataOutW[191:160]; 
assign MEMOCMux17_inw7 = dataOutW[223:192]; 
assign MEMOCMux17_inw8 = dataOutW[255:224]; 
assign MEMOCMux17_inw9 = dataOutW[287:256]; 
assign MEMOCMux17_inw10 = globalDataIn[575:544]; 
assign MEMOCMux17_selw = mOutConfigW[71:68]; 
assign MEMC17_data_out_ctx2 = mDataFromMem[575:544]; 
assign mDataToMem[575:544] = MEMC17_data_in_ctx1; 
assign globalDataOut[575:544] = MEMC17_data_to_Core; 
assign MEMC17_valid_ctx1 = valid1[17:17]; 
assign MEMC17_write_en_ctx1 = WEn1[17:17]; 
assign MEMC17_stride_ctx1 = stride1[17:17]; 
assign MEMC17_start_addr_ctx1 = startAddr1[107:102]; 
assign MEMC17_burst_count_ctx1 = count1[125:119]; 
assign mAddr1[107:102] = MEMC17_addr_out_ctx1; 
assign mEn1[17:17] = MEMC17_mem_en_ctx1; 
assign mWEn1[17:17] = MEMC17_write_mem_en_ctx1; 
assign MEMC17_valid_ctx2 = valid2[17:17]; 
assign MEMC17_write_en_ctx2 = WEn2[17:17]; 
assign MEMC17_stride_ctx2 = stride2[17:17]; 
assign MEMC17_start_addr_ctx2 = startAddr2[107:102]; 
assign mAddr2[107:102] = MEMC17_addr_out_ctx2; 
assign MEMC17_burst_count_ctx2 = count2[125:119]; 
assign mEn2[17:17] = MEMC17_mem_en_ctx2; 
assign mWEn2[17:17] = MEMC17_write_mem_en_ctx2; 
wire [31:0] MEMOCMux18_inw1;
wire [31:0] MEMOCMux18_inw2;
wire [31:0] MEMOCMux18_inw3;
wire [31:0] MEMOCMux18_inw4;
wire [31:0] MEMOCMux18_inw5;
wire [31:0] MEMOCMux18_inw6;
wire [31:0] MEMOCMux18_inw7;
wire [31:0] MEMOCMux18_inw8;
wire [31:0] MEMOCMux18_inw9;
wire [31:0] MEMOCMux18_inw10;
wire [31:0] MEMOCMux18_outw1;
wire [3:0] MEMOCMux18_selw;
HA_10IM MEMOCMux18 (
.DataIn_1(MEMOCMux18_inw1),
.DataIn_2(MEMOCMux18_inw2),
.DataIn_3(MEMOCMux18_inw3),
.DataIn_4(MEMOCMux18_inw4),
.DataIn_5(MEMOCMux18_inw5),
.DataIn_6(MEMOCMux18_inw6),
.DataIn_7(MEMOCMux18_inw7),
.DataIn_8(MEMOCMux18_inw8),
.DataIn_9(MEMOCMux18_inw9),
.DataIn_10(MEMOCMux18_inw10),
.DataOut_1(MEMOCMux18_outw1),
.sel(MEMOCMux18_selw));
defparam MEMOCMux18.Mux_BW = 32;
assign MEMC18_data_from_Core = MEMOCMux18_outw1;
assign MEMOCMux18_inw1 = dataOutW[31:0]; 
assign MEMOCMux18_inw2 = dataOutW[63:32]; 
assign MEMOCMux18_inw3 = dataOutW[95:64]; 
assign MEMOCMux18_inw4 = dataOutW[127:96]; 
assign MEMOCMux18_inw5 = dataOutW[159:128]; 
assign MEMOCMux18_inw6 = dataOutW[191:160]; 
assign MEMOCMux18_inw7 = dataOutW[223:192]; 
assign MEMOCMux18_inw8 = dataOutW[255:224]; 
assign MEMOCMux18_inw9 = dataOutW[287:256]; 
assign MEMOCMux18_inw10 = globalDataIn[607:576]; 
assign MEMOCMux18_selw = mOutConfigW[75:72]; 
assign MEMC18_data_out_ctx2 = mDataFromMem[607:576]; 
assign mDataToMem[607:576] = MEMC18_data_in_ctx1; 
assign globalDataOut[607:576] = MEMC18_data_to_Core; 
assign MEMC18_valid_ctx1 = valid1[18:18]; 
assign MEMC18_write_en_ctx1 = WEn1[18:18]; 
assign MEMC18_stride_ctx1 = stride1[18:18]; 
assign MEMC18_start_addr_ctx1 = startAddr1[113:108]; 
assign MEMC18_burst_count_ctx1 = count1[132:126]; 
assign mAddr1[113:108] = MEMC18_addr_out_ctx1; 
assign mEn1[18:18] = MEMC18_mem_en_ctx1; 
assign mWEn1[18:18] = MEMC18_write_mem_en_ctx1; 
assign MEMC18_valid_ctx2 = valid2[18:18]; 
assign MEMC18_write_en_ctx2 = WEn2[18:18]; 
assign MEMC18_stride_ctx2 = stride2[18:18]; 
assign MEMC18_start_addr_ctx2 = startAddr2[113:108]; 
assign mAddr2[113:108] = MEMC18_addr_out_ctx2; 
assign MEMC18_burst_count_ctx2 = count2[132:126]; 
assign mEn2[18:18] = MEMC18_mem_en_ctx2; 
assign mWEn2[18:18] = MEMC18_write_mem_en_ctx2; 
wire [31:0] MEMOCMux19_inw1;
wire [31:0] MEMOCMux19_inw2;
wire [31:0] MEMOCMux19_inw3;
wire [31:0] MEMOCMux19_inw4;
wire [31:0] MEMOCMux19_inw5;
wire [31:0] MEMOCMux19_inw6;
wire [31:0] MEMOCMux19_inw7;
wire [31:0] MEMOCMux19_inw8;
wire [31:0] MEMOCMux19_inw9;
wire [31:0] MEMOCMux19_inw10;
wire [31:0] MEMOCMux19_outw1;
wire [3:0] MEMOCMux19_selw;
HA_10IM MEMOCMux19 (
.DataIn_1(MEMOCMux19_inw1),
.DataIn_2(MEMOCMux19_inw2),
.DataIn_3(MEMOCMux19_inw3),
.DataIn_4(MEMOCMux19_inw4),
.DataIn_5(MEMOCMux19_inw5),
.DataIn_6(MEMOCMux19_inw6),
.DataIn_7(MEMOCMux19_inw7),
.DataIn_8(MEMOCMux19_inw8),
.DataIn_9(MEMOCMux19_inw9),
.DataIn_10(MEMOCMux19_inw10),
.DataOut_1(MEMOCMux19_outw1),
.sel(MEMOCMux19_selw));
defparam MEMOCMux19.Mux_BW = 32;
assign MEMC19_data_from_Core = MEMOCMux19_outw1;
assign MEMOCMux19_inw1 = dataOutW[31:0]; 
assign MEMOCMux19_inw2 = dataOutW[63:32]; 
assign MEMOCMux19_inw3 = dataOutW[95:64]; 
assign MEMOCMux19_inw4 = dataOutW[127:96]; 
assign MEMOCMux19_inw5 = dataOutW[159:128]; 
assign MEMOCMux19_inw6 = dataOutW[191:160]; 
assign MEMOCMux19_inw7 = dataOutW[223:192]; 
assign MEMOCMux19_inw8 = dataOutW[255:224]; 
assign MEMOCMux19_inw9 = dataOutW[287:256]; 
assign MEMOCMux19_inw10 = globalDataIn[639:608]; 
assign MEMOCMux19_selw = mOutConfigW[79:76]; 
assign MEMC19_data_out_ctx2 = mDataFromMem[639:608]; 
assign mDataToMem[639:608] = MEMC19_data_in_ctx1; 
assign globalDataOut[639:608] = MEMC19_data_to_Core; 
assign MEMC19_valid_ctx1 = valid1[19:19]; 
assign MEMC19_write_en_ctx1 = WEn1[19:19]; 
assign MEMC19_stride_ctx1 = stride1[19:19]; 
assign MEMC19_start_addr_ctx1 = startAddr1[119:114]; 
assign MEMC19_burst_count_ctx1 = count1[139:133]; 
assign mAddr1[119:114] = MEMC19_addr_out_ctx1; 
assign mEn1[19:19] = MEMC19_mem_en_ctx1; 
assign mWEn1[19:19] = MEMC19_write_mem_en_ctx1; 
assign MEMC19_valid_ctx2 = valid2[19:19]; 
assign MEMC19_write_en_ctx2 = WEn2[19:19]; 
assign MEMC19_stride_ctx2 = stride2[19:19]; 
assign MEMC19_start_addr_ctx2 = startAddr2[119:114]; 
assign mAddr2[119:114] = MEMC19_addr_out_ctx2; 
assign MEMC19_burst_count_ctx2 = count2[139:133]; 
assign mEn2[19:19] = MEMC19_mem_en_ctx2; 
assign mWEn2[19:19] = MEMC19_write_mem_en_ctx2; 
wire [31:0] MEMOCMux20_inw1;
wire [31:0] MEMOCMux20_inw2;
wire [31:0] MEMOCMux20_inw3;
wire [31:0] MEMOCMux20_inw4;
wire [31:0] MEMOCMux20_inw5;
wire [31:0] MEMOCMux20_inw6;
wire [31:0] MEMOCMux20_inw7;
wire [31:0] MEMOCMux20_inw8;
wire [31:0] MEMOCMux20_inw9;
wire [31:0] MEMOCMux20_inw10;
wire [31:0] MEMOCMux20_outw1;
wire [3:0] MEMOCMux20_selw;
HA_10IM MEMOCMux20 (
.DataIn_1(MEMOCMux20_inw1),
.DataIn_2(MEMOCMux20_inw2),
.DataIn_3(MEMOCMux20_inw3),
.DataIn_4(MEMOCMux20_inw4),
.DataIn_5(MEMOCMux20_inw5),
.DataIn_6(MEMOCMux20_inw6),
.DataIn_7(MEMOCMux20_inw7),
.DataIn_8(MEMOCMux20_inw8),
.DataIn_9(MEMOCMux20_inw9),
.DataIn_10(MEMOCMux20_inw10),
.DataOut_1(MEMOCMux20_outw1),
.sel(MEMOCMux20_selw));
defparam MEMOCMux20.Mux_BW = 32;
assign MEMC20_data_from_Core = MEMOCMux20_outw1;
assign MEMOCMux20_inw1 = dataOutW[31:0]; 
assign MEMOCMux20_inw2 = dataOutW[63:32]; 
assign MEMOCMux20_inw3 = dataOutW[95:64]; 
assign MEMOCMux20_inw4 = dataOutW[127:96]; 
assign MEMOCMux20_inw5 = dataOutW[159:128]; 
assign MEMOCMux20_inw6 = dataOutW[191:160]; 
assign MEMOCMux20_inw7 = dataOutW[223:192]; 
assign MEMOCMux20_inw8 = dataOutW[255:224]; 
assign MEMOCMux20_inw9 = dataOutW[287:256]; 
assign MEMOCMux20_inw10 = globalDataIn[671:640]; 
assign MEMOCMux20_selw = mOutConfigW[83:80]; 
assign MEMC20_data_out_ctx2 = mDataFromMem[671:640]; 
assign mDataToMem[671:640] = MEMC20_data_in_ctx1; 
assign globalDataOut[671:640] = MEMC20_data_to_Core; 
assign MEMC20_valid_ctx1 = valid1[20:20]; 
assign MEMC20_write_en_ctx1 = WEn1[20:20]; 
assign MEMC20_stride_ctx1 = stride1[20:20]; 
assign MEMC20_start_addr_ctx1 = startAddr1[125:120]; 
assign MEMC20_burst_count_ctx1 = count1[146:140]; 
assign mAddr1[125:120] = MEMC20_addr_out_ctx1; 
assign mEn1[20:20] = MEMC20_mem_en_ctx1; 
assign mWEn1[20:20] = MEMC20_write_mem_en_ctx1; 
assign MEMC20_valid_ctx2 = valid2[20:20]; 
assign MEMC20_write_en_ctx2 = WEn2[20:20]; 
assign MEMC20_stride_ctx2 = stride2[20:20]; 
assign MEMC20_start_addr_ctx2 = startAddr2[125:120]; 
assign mAddr2[125:120] = MEMC20_addr_out_ctx2; 
assign MEMC20_burst_count_ctx2 = count2[146:140]; 
assign mEn2[20:20] = MEMC20_mem_en_ctx2; 
assign mWEn2[20:20] = MEMC20_write_mem_en_ctx2; 
wire [31:0] MEMOCMux21_inw1;
wire [31:0] MEMOCMux21_inw2;
wire [31:0] MEMOCMux21_inw3;
wire [31:0] MEMOCMux21_inw4;
wire [31:0] MEMOCMux21_inw5;
wire [31:0] MEMOCMux21_inw6;
wire [31:0] MEMOCMux21_inw7;
wire [31:0] MEMOCMux21_inw8;
wire [31:0] MEMOCMux21_inw9;
wire [31:0] MEMOCMux21_inw10;
wire [31:0] MEMOCMux21_outw1;
wire [3:0] MEMOCMux21_selw;
HA_10IM MEMOCMux21 (
.DataIn_1(MEMOCMux21_inw1),
.DataIn_2(MEMOCMux21_inw2),
.DataIn_3(MEMOCMux21_inw3),
.DataIn_4(MEMOCMux21_inw4),
.DataIn_5(MEMOCMux21_inw5),
.DataIn_6(MEMOCMux21_inw6),
.DataIn_7(MEMOCMux21_inw7),
.DataIn_8(MEMOCMux21_inw8),
.DataIn_9(MEMOCMux21_inw9),
.DataIn_10(MEMOCMux21_inw10),
.DataOut_1(MEMOCMux21_outw1),
.sel(MEMOCMux21_selw));
defparam MEMOCMux21.Mux_BW = 32;
assign MEMC21_data_from_Core = MEMOCMux21_outw1;
assign MEMOCMux21_inw1 = dataOutW[31:0]; 
assign MEMOCMux21_inw2 = dataOutW[63:32]; 
assign MEMOCMux21_inw3 = dataOutW[95:64]; 
assign MEMOCMux21_inw4 = dataOutW[127:96]; 
assign MEMOCMux21_inw5 = dataOutW[159:128]; 
assign MEMOCMux21_inw6 = dataOutW[191:160]; 
assign MEMOCMux21_inw7 = dataOutW[223:192]; 
assign MEMOCMux21_inw8 = dataOutW[255:224]; 
assign MEMOCMux21_inw9 = dataOutW[287:256]; 
assign MEMOCMux21_inw10 = globalDataIn[703:672]; 
assign MEMOCMux21_selw = mOutConfigW[87:84]; 
assign MEMC21_data_out_ctx2 = mDataFromMem[703:672]; 
assign mDataToMem[703:672] = MEMC21_data_in_ctx1; 
assign globalDataOut[703:672] = MEMC21_data_to_Core; 
assign MEMC21_valid_ctx1 = valid1[21:21]; 
assign MEMC21_write_en_ctx1 = WEn1[21:21]; 
assign MEMC21_stride_ctx1 = stride1[21:21]; 
assign MEMC21_start_addr_ctx1 = startAddr1[131:126]; 
assign MEMC21_burst_count_ctx1 = count1[153:147]; 
assign mAddr1[131:126] = MEMC21_addr_out_ctx1; 
assign mEn1[21:21] = MEMC21_mem_en_ctx1; 
assign mWEn1[21:21] = MEMC21_write_mem_en_ctx1; 
assign MEMC21_valid_ctx2 = valid2[21:21]; 
assign MEMC21_write_en_ctx2 = WEn2[21:21]; 
assign MEMC21_stride_ctx2 = stride2[21:21]; 
assign MEMC21_start_addr_ctx2 = startAddr2[131:126]; 
assign mAddr2[131:126] = MEMC21_addr_out_ctx2; 
assign MEMC21_burst_count_ctx2 = count2[153:147]; 
assign mEn2[21:21] = MEMC21_mem_en_ctx2; 
assign mWEn2[21:21] = MEMC21_write_mem_en_ctx2; 
wire [31:0] MEMOCMux22_inw1;
wire [31:0] MEMOCMux22_inw2;
wire [31:0] MEMOCMux22_inw3;
wire [31:0] MEMOCMux22_inw4;
wire [31:0] MEMOCMux22_inw5;
wire [31:0] MEMOCMux22_inw6;
wire [31:0] MEMOCMux22_inw7;
wire [31:0] MEMOCMux22_inw8;
wire [31:0] MEMOCMux22_inw9;
wire [31:0] MEMOCMux22_inw10;
wire [31:0] MEMOCMux22_outw1;
wire [3:0] MEMOCMux22_selw;
HA_10IM MEMOCMux22 (
.DataIn_1(MEMOCMux22_inw1),
.DataIn_2(MEMOCMux22_inw2),
.DataIn_3(MEMOCMux22_inw3),
.DataIn_4(MEMOCMux22_inw4),
.DataIn_5(MEMOCMux22_inw5),
.DataIn_6(MEMOCMux22_inw6),
.DataIn_7(MEMOCMux22_inw7),
.DataIn_8(MEMOCMux22_inw8),
.DataIn_9(MEMOCMux22_inw9),
.DataIn_10(MEMOCMux22_inw10),
.DataOut_1(MEMOCMux22_outw1),
.sel(MEMOCMux22_selw));
defparam MEMOCMux22.Mux_BW = 32;
assign MEMC22_data_from_Core = MEMOCMux22_outw1;
assign MEMOCMux22_inw1 = dataOutW[31:0]; 
assign MEMOCMux22_inw2 = dataOutW[63:32]; 
assign MEMOCMux22_inw3 = dataOutW[95:64]; 
assign MEMOCMux22_inw4 = dataOutW[127:96]; 
assign MEMOCMux22_inw5 = dataOutW[159:128]; 
assign MEMOCMux22_inw6 = dataOutW[191:160]; 
assign MEMOCMux22_inw7 = dataOutW[223:192]; 
assign MEMOCMux22_inw8 = dataOutW[255:224]; 
assign MEMOCMux22_inw9 = dataOutW[287:256]; 
assign MEMOCMux22_inw10 = globalDataIn[735:704]; 
assign MEMOCMux22_selw = mOutConfigW[91:88]; 
assign MEMC22_data_out_ctx2 = mDataFromMem[735:704]; 
assign mDataToMem[735:704] = MEMC22_data_in_ctx1; 
assign globalDataOut[735:704] = MEMC22_data_to_Core; 
assign MEMC22_valid_ctx1 = valid1[22:22]; 
assign MEMC22_write_en_ctx1 = WEn1[22:22]; 
assign MEMC22_stride_ctx1 = stride1[22:22]; 
assign MEMC22_start_addr_ctx1 = startAddr1[137:132]; 
assign MEMC22_burst_count_ctx1 = count1[160:154]; 
assign mAddr1[137:132] = MEMC22_addr_out_ctx1; 
assign mEn1[22:22] = MEMC22_mem_en_ctx1; 
assign mWEn1[22:22] = MEMC22_write_mem_en_ctx1; 
assign MEMC22_valid_ctx2 = valid2[22:22]; 
assign MEMC22_write_en_ctx2 = WEn2[22:22]; 
assign MEMC22_stride_ctx2 = stride2[22:22]; 
assign MEMC22_start_addr_ctx2 = startAddr2[137:132]; 
assign mAddr2[137:132] = MEMC22_addr_out_ctx2; 
assign MEMC22_burst_count_ctx2 = count2[160:154]; 
assign mEn2[22:22] = MEMC22_mem_en_ctx2; 
assign mWEn2[22:22] = MEMC22_write_mem_en_ctx2; 
wire [31:0] MEMOCMux23_inw1;
wire [31:0] MEMOCMux23_inw2;
wire [31:0] MEMOCMux23_inw3;
wire [31:0] MEMOCMux23_inw4;
wire [31:0] MEMOCMux23_inw5;
wire [31:0] MEMOCMux23_inw6;
wire [31:0] MEMOCMux23_inw7;
wire [31:0] MEMOCMux23_inw8;
wire [31:0] MEMOCMux23_inw9;
wire [31:0] MEMOCMux23_inw10;
wire [31:0] MEMOCMux23_outw1;
wire [3:0] MEMOCMux23_selw;
HA_10IM MEMOCMux23 (
.DataIn_1(MEMOCMux23_inw1),
.DataIn_2(MEMOCMux23_inw2),
.DataIn_3(MEMOCMux23_inw3),
.DataIn_4(MEMOCMux23_inw4),
.DataIn_5(MEMOCMux23_inw5),
.DataIn_6(MEMOCMux23_inw6),
.DataIn_7(MEMOCMux23_inw7),
.DataIn_8(MEMOCMux23_inw8),
.DataIn_9(MEMOCMux23_inw9),
.DataIn_10(MEMOCMux23_inw10),
.DataOut_1(MEMOCMux23_outw1),
.sel(MEMOCMux23_selw));
defparam MEMOCMux23.Mux_BW = 32;
assign MEMC23_data_from_Core = MEMOCMux23_outw1;
assign MEMOCMux23_inw1 = dataOutW[31:0]; 
assign MEMOCMux23_inw2 = dataOutW[63:32]; 
assign MEMOCMux23_inw3 = dataOutW[95:64]; 
assign MEMOCMux23_inw4 = dataOutW[127:96]; 
assign MEMOCMux23_inw5 = dataOutW[159:128]; 
assign MEMOCMux23_inw6 = dataOutW[191:160]; 
assign MEMOCMux23_inw7 = dataOutW[223:192]; 
assign MEMOCMux23_inw8 = dataOutW[255:224]; 
assign MEMOCMux23_inw9 = dataOutW[287:256]; 
assign MEMOCMux23_inw10 = globalDataIn[767:736]; 
assign MEMOCMux23_selw = mOutConfigW[95:92]; 
assign MEMC23_data_out_ctx2 = mDataFromMem[767:736]; 
assign mDataToMem[767:736] = MEMC23_data_in_ctx1; 
assign globalDataOut[767:736] = MEMC23_data_to_Core; 
assign MEMC23_valid_ctx1 = valid1[23:23]; 
assign MEMC23_write_en_ctx1 = WEn1[23:23]; 
assign MEMC23_stride_ctx1 = stride1[23:23]; 
assign MEMC23_start_addr_ctx1 = startAddr1[143:138]; 
assign MEMC23_burst_count_ctx1 = count1[167:161]; 
assign mAddr1[143:138] = MEMC23_addr_out_ctx1; 
assign mEn1[23:23] = MEMC23_mem_en_ctx1; 
assign mWEn1[23:23] = MEMC23_write_mem_en_ctx1; 
assign MEMC23_valid_ctx2 = valid2[23:23]; 
assign MEMC23_write_en_ctx2 = WEn2[23:23]; 
assign MEMC23_stride_ctx2 = stride2[23:23]; 
assign MEMC23_start_addr_ctx2 = startAddr2[143:138]; 
assign mAddr2[143:138] = MEMC23_addr_out_ctx2; 
assign MEMC23_burst_count_ctx2 = count2[167:161]; 
assign mEn2[23:23] = MEMC23_mem_en_ctx2; 
assign mWEn2[23:23] = MEMC23_write_mem_en_ctx2; 
wire [31:0] MEMOCMux24_inw1;
wire [31:0] MEMOCMux24_inw2;
wire [31:0] MEMOCMux24_inw3;
wire [31:0] MEMOCMux24_inw4;
wire [31:0] MEMOCMux24_inw5;
wire [31:0] MEMOCMux24_inw6;
wire [31:0] MEMOCMux24_inw7;
wire [31:0] MEMOCMux24_inw8;
wire [31:0] MEMOCMux24_inw9;
wire [31:0] MEMOCMux24_inw10;
wire [31:0] MEMOCMux24_outw1;
wire [3:0] MEMOCMux24_selw;
HA_10IM MEMOCMux24 (
.DataIn_1(MEMOCMux24_inw1),
.DataIn_2(MEMOCMux24_inw2),
.DataIn_3(MEMOCMux24_inw3),
.DataIn_4(MEMOCMux24_inw4),
.DataIn_5(MEMOCMux24_inw5),
.DataIn_6(MEMOCMux24_inw6),
.DataIn_7(MEMOCMux24_inw7),
.DataIn_8(MEMOCMux24_inw8),
.DataIn_9(MEMOCMux24_inw9),
.DataIn_10(MEMOCMux24_inw10),
.DataOut_1(MEMOCMux24_outw1),
.sel(MEMOCMux24_selw));
defparam MEMOCMux24.Mux_BW = 32;
assign MEMC24_data_from_Core = MEMOCMux24_outw1;
assign MEMOCMux24_inw1 = dataOutW[31:0]; 
assign MEMOCMux24_inw2 = dataOutW[63:32]; 
assign MEMOCMux24_inw3 = dataOutW[95:64]; 
assign MEMOCMux24_inw4 = dataOutW[127:96]; 
assign MEMOCMux24_inw5 = dataOutW[159:128]; 
assign MEMOCMux24_inw6 = dataOutW[191:160]; 
assign MEMOCMux24_inw7 = dataOutW[223:192]; 
assign MEMOCMux24_inw8 = dataOutW[255:224]; 
assign MEMOCMux24_inw9 = dataOutW[287:256]; 
assign MEMOCMux24_inw10 = globalDataIn[799:768]; 
assign MEMOCMux24_selw = mOutConfigW[99:96]; 
assign MEMC24_data_out_ctx2 = mDataFromMem[799:768]; 
assign mDataToMem[799:768] = MEMC24_data_in_ctx1; 
assign globalDataOut[799:768] = MEMC24_data_to_Core; 
assign MEMC24_valid_ctx1 = valid1[24:24]; 
assign MEMC24_write_en_ctx1 = WEn1[24:24]; 
assign MEMC24_stride_ctx1 = stride1[24:24]; 
assign MEMC24_start_addr_ctx1 = startAddr1[149:144]; 
assign MEMC24_burst_count_ctx1 = count1[174:168]; 
assign mAddr1[149:144] = MEMC24_addr_out_ctx1; 
assign mEn1[24:24] = MEMC24_mem_en_ctx1; 
assign mWEn1[24:24] = MEMC24_write_mem_en_ctx1; 
assign MEMC24_valid_ctx2 = valid2[24:24]; 
assign MEMC24_write_en_ctx2 = WEn2[24:24]; 
assign MEMC24_stride_ctx2 = stride2[24:24]; 
assign MEMC24_start_addr_ctx2 = startAddr2[149:144]; 
assign mAddr2[149:144] = MEMC24_addr_out_ctx2; 
assign MEMC24_burst_count_ctx2 = count2[174:168]; 
assign mEn2[24:24] = MEMC24_mem_en_ctx2; 
assign mWEn2[24:24] = MEMC24_write_mem_en_ctx2; 
wire [31:0] MEMOCMux25_inw1;
wire [31:0] MEMOCMux25_inw2;
wire [31:0] MEMOCMux25_inw3;
wire [31:0] MEMOCMux25_inw4;
wire [31:0] MEMOCMux25_inw5;
wire [31:0] MEMOCMux25_inw6;
wire [31:0] MEMOCMux25_inw7;
wire [31:0] MEMOCMux25_inw8;
wire [31:0] MEMOCMux25_inw9;
wire [31:0] MEMOCMux25_inw10;
wire [31:0] MEMOCMux25_outw1;
wire [3:0] MEMOCMux25_selw;
HA_10IM MEMOCMux25 (
.DataIn_1(MEMOCMux25_inw1),
.DataIn_2(MEMOCMux25_inw2),
.DataIn_3(MEMOCMux25_inw3),
.DataIn_4(MEMOCMux25_inw4),
.DataIn_5(MEMOCMux25_inw5),
.DataIn_6(MEMOCMux25_inw6),
.DataIn_7(MEMOCMux25_inw7),
.DataIn_8(MEMOCMux25_inw8),
.DataIn_9(MEMOCMux25_inw9),
.DataIn_10(MEMOCMux25_inw10),
.DataOut_1(MEMOCMux25_outw1),
.sel(MEMOCMux25_selw));
defparam MEMOCMux25.Mux_BW = 32;
assign MEMC25_data_from_Core = MEMOCMux25_outw1;
assign MEMOCMux25_inw1 = dataOutW[31:0]; 
assign MEMOCMux25_inw2 = dataOutW[63:32]; 
assign MEMOCMux25_inw3 = dataOutW[95:64]; 
assign MEMOCMux25_inw4 = dataOutW[127:96]; 
assign MEMOCMux25_inw5 = dataOutW[159:128]; 
assign MEMOCMux25_inw6 = dataOutW[191:160]; 
assign MEMOCMux25_inw7 = dataOutW[223:192]; 
assign MEMOCMux25_inw8 = dataOutW[255:224]; 
assign MEMOCMux25_inw9 = dataOutW[287:256]; 
assign MEMOCMux25_inw10 = globalDataIn[831:800]; 
assign MEMOCMux25_selw = mOutConfigW[103:100]; 
assign MEMC25_data_out_ctx2 = mDataFromMem[831:800]; 
assign mDataToMem[831:800] = MEMC25_data_in_ctx1; 
assign globalDataOut[831:800] = MEMC25_data_to_Core; 
assign MEMC25_valid_ctx1 = valid1[25:25]; 
assign MEMC25_write_en_ctx1 = WEn1[25:25]; 
assign MEMC25_stride_ctx1 = stride1[25:25]; 
assign MEMC25_start_addr_ctx1 = startAddr1[155:150]; 
assign MEMC25_burst_count_ctx1 = count1[181:175]; 
assign mAddr1[155:150] = MEMC25_addr_out_ctx1; 
assign mEn1[25:25] = MEMC25_mem_en_ctx1; 
assign mWEn1[25:25] = MEMC25_write_mem_en_ctx1; 
assign MEMC25_valid_ctx2 = valid2[25:25]; 
assign MEMC25_write_en_ctx2 = WEn2[25:25]; 
assign MEMC25_stride_ctx2 = stride2[25:25]; 
assign MEMC25_start_addr_ctx2 = startAddr2[155:150]; 
assign mAddr2[155:150] = MEMC25_addr_out_ctx2; 
assign MEMC25_burst_count_ctx2 = count2[181:175]; 
assign mEn2[25:25] = MEMC25_mem_en_ctx2; 
assign mWEn2[25:25] = MEMC25_write_mem_en_ctx2; 
wire [31:0] MEMOCMux26_inw1;
wire [31:0] MEMOCMux26_inw2;
wire [31:0] MEMOCMux26_inw3;
wire [31:0] MEMOCMux26_inw4;
wire [31:0] MEMOCMux26_inw5;
wire [31:0] MEMOCMux26_inw6;
wire [31:0] MEMOCMux26_inw7;
wire [31:0] MEMOCMux26_inw8;
wire [31:0] MEMOCMux26_inw9;
wire [31:0] MEMOCMux26_inw10;
wire [31:0] MEMOCMux26_outw1;
wire [3:0] MEMOCMux26_selw;
HA_10IM MEMOCMux26 (
.DataIn_1(MEMOCMux26_inw1),
.DataIn_2(MEMOCMux26_inw2),
.DataIn_3(MEMOCMux26_inw3),
.DataIn_4(MEMOCMux26_inw4),
.DataIn_5(MEMOCMux26_inw5),
.DataIn_6(MEMOCMux26_inw6),
.DataIn_7(MEMOCMux26_inw7),
.DataIn_8(MEMOCMux26_inw8),
.DataIn_9(MEMOCMux26_inw9),
.DataIn_10(MEMOCMux26_inw10),
.DataOut_1(MEMOCMux26_outw1),
.sel(MEMOCMux26_selw));
defparam MEMOCMux26.Mux_BW = 32;
assign MEMC26_data_from_Core = MEMOCMux26_outw1;
assign MEMOCMux26_inw1 = dataOutW[31:0]; 
assign MEMOCMux26_inw2 = dataOutW[63:32]; 
assign MEMOCMux26_inw3 = dataOutW[95:64]; 
assign MEMOCMux26_inw4 = dataOutW[127:96]; 
assign MEMOCMux26_inw5 = dataOutW[159:128]; 
assign MEMOCMux26_inw6 = dataOutW[191:160]; 
assign MEMOCMux26_inw7 = dataOutW[223:192]; 
assign MEMOCMux26_inw8 = dataOutW[255:224]; 
assign MEMOCMux26_inw9 = dataOutW[287:256]; 
assign MEMOCMux26_inw10 = globalDataIn[863:832]; 
assign MEMOCMux26_selw = mOutConfigW[107:104]; 
assign MEMC26_data_out_ctx2 = mDataFromMem[863:832]; 
assign mDataToMem[863:832] = MEMC26_data_in_ctx1; 
assign globalDataOut[863:832] = MEMC26_data_to_Core; 
assign MEMC26_valid_ctx1 = valid1[26:26]; 
assign MEMC26_write_en_ctx1 = WEn1[26:26]; 
assign MEMC26_stride_ctx1 = stride1[26:26]; 
assign MEMC26_start_addr_ctx1 = startAddr1[161:156]; 
assign MEMC26_burst_count_ctx1 = count1[188:182]; 
assign mAddr1[161:156] = MEMC26_addr_out_ctx1; 
assign mEn1[26:26] = MEMC26_mem_en_ctx1; 
assign mWEn1[26:26] = MEMC26_write_mem_en_ctx1; 
assign MEMC26_valid_ctx2 = valid2[26:26]; 
assign MEMC26_write_en_ctx2 = WEn2[26:26]; 
assign MEMC26_stride_ctx2 = stride2[26:26]; 
assign MEMC26_start_addr_ctx2 = startAddr2[161:156]; 
assign mAddr2[161:156] = MEMC26_addr_out_ctx2; 
assign MEMC26_burst_count_ctx2 = count2[188:182]; 
assign mEn2[26:26] = MEMC26_mem_en_ctx2; 
assign mWEn2[26:26] = MEMC26_write_mem_en_ctx2; 
wire [31:0] MEMOCMux27_inw1;
wire [31:0] MEMOCMux27_inw2;
wire [31:0] MEMOCMux27_inw3;
wire [31:0] MEMOCMux27_inw4;
wire [31:0] MEMOCMux27_inw5;
wire [31:0] MEMOCMux27_inw6;
wire [31:0] MEMOCMux27_inw7;
wire [31:0] MEMOCMux27_inw8;
wire [31:0] MEMOCMux27_inw9;
wire [31:0] MEMOCMux27_inw10;
wire [31:0] MEMOCMux27_outw1;
wire [3:0] MEMOCMux27_selw;
HA_10IM MEMOCMux27 (
.DataIn_1(MEMOCMux27_inw1),
.DataIn_2(MEMOCMux27_inw2),
.DataIn_3(MEMOCMux27_inw3),
.DataIn_4(MEMOCMux27_inw4),
.DataIn_5(MEMOCMux27_inw5),
.DataIn_6(MEMOCMux27_inw6),
.DataIn_7(MEMOCMux27_inw7),
.DataIn_8(MEMOCMux27_inw8),
.DataIn_9(MEMOCMux27_inw9),
.DataIn_10(MEMOCMux27_inw10),
.DataOut_1(MEMOCMux27_outw1),
.sel(MEMOCMux27_selw));
defparam MEMOCMux27.Mux_BW = 32;
assign MEMC27_data_from_Core = MEMOCMux27_outw1;
assign MEMOCMux27_inw1 = dataOutW[31:0]; 
assign MEMOCMux27_inw2 = dataOutW[63:32]; 
assign MEMOCMux27_inw3 = dataOutW[95:64]; 
assign MEMOCMux27_inw4 = dataOutW[127:96]; 
assign MEMOCMux27_inw5 = dataOutW[159:128]; 
assign MEMOCMux27_inw6 = dataOutW[191:160]; 
assign MEMOCMux27_inw7 = dataOutW[223:192]; 
assign MEMOCMux27_inw8 = dataOutW[255:224]; 
assign MEMOCMux27_inw9 = dataOutW[287:256]; 
assign MEMOCMux27_inw10 = globalDataIn[895:864]; 
assign MEMOCMux27_selw = mOutConfigW[111:108]; 
assign MEMC27_data_out_ctx2 = mDataFromMem[895:864]; 
assign mDataToMem[895:864] = MEMC27_data_in_ctx1; 
assign globalDataOut[895:864] = MEMC27_data_to_Core; 
assign MEMC27_valid_ctx1 = valid1[27:27]; 
assign MEMC27_write_en_ctx1 = WEn1[27:27]; 
assign MEMC27_stride_ctx1 = stride1[27:27]; 
assign MEMC27_start_addr_ctx1 = startAddr1[167:162]; 
assign MEMC27_burst_count_ctx1 = count1[195:189]; 
assign mAddr1[167:162] = MEMC27_addr_out_ctx1; 
assign mEn1[27:27] = MEMC27_mem_en_ctx1; 
assign mWEn1[27:27] = MEMC27_write_mem_en_ctx1; 
assign MEMC27_valid_ctx2 = valid2[27:27]; 
assign MEMC27_write_en_ctx2 = WEn2[27:27]; 
assign MEMC27_stride_ctx2 = stride2[27:27]; 
assign MEMC27_start_addr_ctx2 = startAddr2[167:162]; 
assign mAddr2[167:162] = MEMC27_addr_out_ctx2; 
assign MEMC27_burst_count_ctx2 = count2[195:189]; 
assign mEn2[27:27] = MEMC27_mem_en_ctx2; 
assign mWEn2[27:27] = MEMC27_write_mem_en_ctx2; 
wire [31:0] MEMOCMux28_inw1;
wire [31:0] MEMOCMux28_inw2;
wire [31:0] MEMOCMux28_inw3;
wire [31:0] MEMOCMux28_inw4;
wire [31:0] MEMOCMux28_inw5;
wire [31:0] MEMOCMux28_inw6;
wire [31:0] MEMOCMux28_inw7;
wire [31:0] MEMOCMux28_inw8;
wire [31:0] MEMOCMux28_inw9;
wire [31:0] MEMOCMux28_inw10;
wire [31:0] MEMOCMux28_outw1;
wire [3:0] MEMOCMux28_selw;
HA_10IM MEMOCMux28 (
.DataIn_1(MEMOCMux28_inw1),
.DataIn_2(MEMOCMux28_inw2),
.DataIn_3(MEMOCMux28_inw3),
.DataIn_4(MEMOCMux28_inw4),
.DataIn_5(MEMOCMux28_inw5),
.DataIn_6(MEMOCMux28_inw6),
.DataIn_7(MEMOCMux28_inw7),
.DataIn_8(MEMOCMux28_inw8),
.DataIn_9(MEMOCMux28_inw9),
.DataIn_10(MEMOCMux28_inw10),
.DataOut_1(MEMOCMux28_outw1),
.sel(MEMOCMux28_selw));
defparam MEMOCMux28.Mux_BW = 32;
assign MEMC28_data_from_Core = MEMOCMux28_outw1;
assign MEMOCMux28_inw1 = dataOutW[31:0]; 
assign MEMOCMux28_inw2 = dataOutW[63:32]; 
assign MEMOCMux28_inw3 = dataOutW[95:64]; 
assign MEMOCMux28_inw4 = dataOutW[127:96]; 
assign MEMOCMux28_inw5 = dataOutW[159:128]; 
assign MEMOCMux28_inw6 = dataOutW[191:160]; 
assign MEMOCMux28_inw7 = dataOutW[223:192]; 
assign MEMOCMux28_inw8 = dataOutW[255:224]; 
assign MEMOCMux28_inw9 = dataOutW[287:256]; 
assign MEMOCMux28_inw10 = globalDataIn[927:896]; 
assign MEMOCMux28_selw = mOutConfigW[115:112]; 
assign MEMC28_data_out_ctx2 = mDataFromMem[927:896]; 
assign mDataToMem[927:896] = MEMC28_data_in_ctx1; 
assign globalDataOut[927:896] = MEMC28_data_to_Core; 
assign MEMC28_valid_ctx1 = valid1[28:28]; 
assign MEMC28_write_en_ctx1 = WEn1[28:28]; 
assign MEMC28_stride_ctx1 = stride1[28:28]; 
assign MEMC28_start_addr_ctx1 = startAddr1[173:168]; 
assign MEMC28_burst_count_ctx1 = count1[202:196]; 
assign mAddr1[173:168] = MEMC28_addr_out_ctx1; 
assign mEn1[28:28] = MEMC28_mem_en_ctx1; 
assign mWEn1[28:28] = MEMC28_write_mem_en_ctx1; 
assign MEMC28_valid_ctx2 = valid2[28:28]; 
assign MEMC28_write_en_ctx2 = WEn2[28:28]; 
assign MEMC28_stride_ctx2 = stride2[28:28]; 
assign MEMC28_start_addr_ctx2 = startAddr2[173:168]; 
assign mAddr2[173:168] = MEMC28_addr_out_ctx2; 
assign MEMC28_burst_count_ctx2 = count2[202:196]; 
assign mEn2[28:28] = MEMC28_mem_en_ctx2; 
assign mWEn2[28:28] = MEMC28_write_mem_en_ctx2; 
wire [31:0] MEMOCMux29_inw1;
wire [31:0] MEMOCMux29_inw2;
wire [31:0] MEMOCMux29_inw3;
wire [31:0] MEMOCMux29_inw4;
wire [31:0] MEMOCMux29_inw5;
wire [31:0] MEMOCMux29_inw6;
wire [31:0] MEMOCMux29_inw7;
wire [31:0] MEMOCMux29_inw8;
wire [31:0] MEMOCMux29_inw9;
wire [31:0] MEMOCMux29_inw10;
wire [31:0] MEMOCMux29_outw1;
wire [3:0] MEMOCMux29_selw;
HA_10IM MEMOCMux29 (
.DataIn_1(MEMOCMux29_inw1),
.DataIn_2(MEMOCMux29_inw2),
.DataIn_3(MEMOCMux29_inw3),
.DataIn_4(MEMOCMux29_inw4),
.DataIn_5(MEMOCMux29_inw5),
.DataIn_6(MEMOCMux29_inw6),
.DataIn_7(MEMOCMux29_inw7),
.DataIn_8(MEMOCMux29_inw8),
.DataIn_9(MEMOCMux29_inw9),
.DataIn_10(MEMOCMux29_inw10),
.DataOut_1(MEMOCMux29_outw1),
.sel(MEMOCMux29_selw));
defparam MEMOCMux29.Mux_BW = 32;
assign MEMC29_data_from_Core = MEMOCMux29_outw1;
assign MEMOCMux29_inw1 = dataOutW[31:0]; 
assign MEMOCMux29_inw2 = dataOutW[63:32]; 
assign MEMOCMux29_inw3 = dataOutW[95:64]; 
assign MEMOCMux29_inw4 = dataOutW[127:96]; 
assign MEMOCMux29_inw5 = dataOutW[159:128]; 
assign MEMOCMux29_inw6 = dataOutW[191:160]; 
assign MEMOCMux29_inw7 = dataOutW[223:192]; 
assign MEMOCMux29_inw8 = dataOutW[255:224]; 
assign MEMOCMux29_inw9 = dataOutW[287:256]; 
assign MEMOCMux29_inw10 = globalDataIn[959:928]; 
assign MEMOCMux29_selw = mOutConfigW[119:116]; 
assign MEMC29_data_out_ctx2 = mDataFromMem[959:928]; 
assign mDataToMem[959:928] = MEMC29_data_in_ctx1; 
assign globalDataOut[959:928] = MEMC29_data_to_Core; 
assign MEMC29_valid_ctx1 = valid1[29:29]; 
assign MEMC29_write_en_ctx1 = WEn1[29:29]; 
assign MEMC29_stride_ctx1 = stride1[29:29]; 
assign MEMC29_start_addr_ctx1 = startAddr1[179:174]; 
assign MEMC29_burst_count_ctx1 = count1[209:203]; 
assign mAddr1[179:174] = MEMC29_addr_out_ctx1; 
assign mEn1[29:29] = MEMC29_mem_en_ctx1; 
assign mWEn1[29:29] = MEMC29_write_mem_en_ctx1; 
assign MEMC29_valid_ctx2 = valid2[29:29]; 
assign MEMC29_write_en_ctx2 = WEn2[29:29]; 
assign MEMC29_stride_ctx2 = stride2[29:29]; 
assign MEMC29_start_addr_ctx2 = startAddr2[179:174]; 
assign mAddr2[179:174] = MEMC29_addr_out_ctx2; 
assign MEMC29_burst_count_ctx2 = count2[209:203]; 
assign mEn2[29:29] = MEMC29_mem_en_ctx2; 
assign mWEn2[29:29] = MEMC29_write_mem_en_ctx2; 
wire [31:0] MEMOCMux30_inw1;
wire [31:0] MEMOCMux30_inw2;
wire [31:0] MEMOCMux30_inw3;
wire [31:0] MEMOCMux30_inw4;
wire [31:0] MEMOCMux30_inw5;
wire [31:0] MEMOCMux30_inw6;
wire [31:0] MEMOCMux30_inw7;
wire [31:0] MEMOCMux30_inw8;
wire [31:0] MEMOCMux30_inw9;
wire [31:0] MEMOCMux30_inw10;
wire [31:0] MEMOCMux30_outw1;
wire [3:0] MEMOCMux30_selw;
HA_10IM MEMOCMux30 (
.DataIn_1(MEMOCMux30_inw1),
.DataIn_2(MEMOCMux30_inw2),
.DataIn_3(MEMOCMux30_inw3),
.DataIn_4(MEMOCMux30_inw4),
.DataIn_5(MEMOCMux30_inw5),
.DataIn_6(MEMOCMux30_inw6),
.DataIn_7(MEMOCMux30_inw7),
.DataIn_8(MEMOCMux30_inw8),
.DataIn_9(MEMOCMux30_inw9),
.DataIn_10(MEMOCMux30_inw10),
.DataOut_1(MEMOCMux30_outw1),
.sel(MEMOCMux30_selw));
defparam MEMOCMux30.Mux_BW = 32;
assign MEMC30_data_from_Core = MEMOCMux30_outw1;
assign MEMOCMux30_inw1 = dataOutW[31:0]; 
assign MEMOCMux30_inw2 = dataOutW[63:32]; 
assign MEMOCMux30_inw3 = dataOutW[95:64]; 
assign MEMOCMux30_inw4 = dataOutW[127:96]; 
assign MEMOCMux30_inw5 = dataOutW[159:128]; 
assign MEMOCMux30_inw6 = dataOutW[191:160]; 
assign MEMOCMux30_inw7 = dataOutW[223:192]; 
assign MEMOCMux30_inw8 = dataOutW[255:224]; 
assign MEMOCMux30_inw9 = dataOutW[287:256]; 
assign MEMOCMux30_inw10 = globalDataIn[991:960]; 
assign MEMOCMux30_selw = mOutConfigW[123:120]; 
assign MEMC30_data_out_ctx2 = mDataFromMem[991:960]; 
assign mDataToMem[991:960] = MEMC30_data_in_ctx1; 
assign globalDataOut[991:960] = MEMC30_data_to_Core; 
assign MEMC30_valid_ctx1 = valid1[30:30]; 
assign MEMC30_write_en_ctx1 = WEn1[30:30]; 
assign MEMC30_stride_ctx1 = stride1[30:30]; 
assign MEMC30_start_addr_ctx1 = startAddr1[185:180]; 
assign MEMC30_burst_count_ctx1 = count1[216:210]; 
assign mAddr1[185:180] = MEMC30_addr_out_ctx1; 
assign mEn1[30:30] = MEMC30_mem_en_ctx1; 
assign mWEn1[30:30] = MEMC30_write_mem_en_ctx1; 
assign MEMC30_valid_ctx2 = valid2[30:30]; 
assign MEMC30_write_en_ctx2 = WEn2[30:30]; 
assign MEMC30_stride_ctx2 = stride2[30:30]; 
assign MEMC30_start_addr_ctx2 = startAddr2[185:180]; 
assign mAddr2[185:180] = MEMC30_addr_out_ctx2; 
assign MEMC30_burst_count_ctx2 = count2[216:210]; 
assign mEn2[30:30] = MEMC30_mem_en_ctx2; 
assign mWEn2[30:30] = MEMC30_write_mem_en_ctx2; 
wire [31:0] MEMOCMux31_inw1;
wire [31:0] MEMOCMux31_inw2;
wire [31:0] MEMOCMux31_inw3;
wire [31:0] MEMOCMux31_inw4;
wire [31:0] MEMOCMux31_inw5;
wire [31:0] MEMOCMux31_inw6;
wire [31:0] MEMOCMux31_inw7;
wire [31:0] MEMOCMux31_inw8;
wire [31:0] MEMOCMux31_inw9;
wire [31:0] MEMOCMux31_inw10;
wire [31:0] MEMOCMux31_outw1;
wire [3:0] MEMOCMux31_selw;
HA_10IM MEMOCMux31 (
.DataIn_1(MEMOCMux31_inw1),
.DataIn_2(MEMOCMux31_inw2),
.DataIn_3(MEMOCMux31_inw3),
.DataIn_4(MEMOCMux31_inw4),
.DataIn_5(MEMOCMux31_inw5),
.DataIn_6(MEMOCMux31_inw6),
.DataIn_7(MEMOCMux31_inw7),
.DataIn_8(MEMOCMux31_inw8),
.DataIn_9(MEMOCMux31_inw9),
.DataIn_10(MEMOCMux31_inw10),
.DataOut_1(MEMOCMux31_outw1),
.sel(MEMOCMux31_selw));
defparam MEMOCMux31.Mux_BW = 32;
assign MEMC31_data_from_Core = MEMOCMux31_outw1;
assign MEMOCMux31_inw1 = dataOutW[31:0]; 
assign MEMOCMux31_inw2 = dataOutW[63:32]; 
assign MEMOCMux31_inw3 = dataOutW[95:64]; 
assign MEMOCMux31_inw4 = dataOutW[127:96]; 
assign MEMOCMux31_inw5 = dataOutW[159:128]; 
assign MEMOCMux31_inw6 = dataOutW[191:160]; 
assign MEMOCMux31_inw7 = dataOutW[223:192]; 
assign MEMOCMux31_inw8 = dataOutW[255:224]; 
assign MEMOCMux31_inw9 = dataOutW[287:256]; 
assign MEMOCMux31_inw10 = globalDataIn[1023:992]; 
assign MEMOCMux31_selw = mOutConfigW[127:124]; 
assign MEMC31_data_out_ctx2 = mDataFromMem[1023:992]; 
assign mDataToMem[1023:992] = MEMC31_data_in_ctx1; 
assign globalDataOut[1023:992] = MEMC31_data_to_Core; 
assign MEMC31_valid_ctx1 = valid1[31:31]; 
assign MEMC31_write_en_ctx1 = WEn1[31:31]; 
assign MEMC31_stride_ctx1 = stride1[31:31]; 
assign MEMC31_start_addr_ctx1 = startAddr1[191:186]; 
assign MEMC31_burst_count_ctx1 = count1[223:217]; 
assign mAddr1[191:186] = MEMC31_addr_out_ctx1; 
assign mEn1[31:31] = MEMC31_mem_en_ctx1; 
assign mWEn1[31:31] = MEMC31_write_mem_en_ctx1; 
assign MEMC31_valid_ctx2 = valid2[31:31]; 
assign MEMC31_write_en_ctx2 = WEn2[31:31]; 
assign MEMC31_stride_ctx2 = stride2[31:31]; 
assign MEMC31_start_addr_ctx2 = startAddr2[191:186]; 
assign mAddr2[191:186] = MEMC31_addr_out_ctx2; 
assign MEMC31_burst_count_ctx2 = count2[223:217]; 
assign mEn2[31:31] = MEMC31_mem_en_ctx2; 
assign mWEn2[31:31] = MEMC31_write_mem_en_ctx2; 
wire [31:0] MEMOCMux32_inw1;
wire [31:0] MEMOCMux32_inw2;
wire [31:0] MEMOCMux32_inw3;
wire [31:0] MEMOCMux32_inw4;
wire [31:0] MEMOCMux32_inw5;
wire [31:0] MEMOCMux32_inw6;
wire [31:0] MEMOCMux32_inw7;
wire [31:0] MEMOCMux32_inw8;
wire [31:0] MEMOCMux32_inw9;
wire [31:0] MEMOCMux32_inw10;
wire [31:0] MEMOCMux32_outw1;
wire [3:0] MEMOCMux32_selw;
HA_10IM MEMOCMux32 (
.DataIn_1(MEMOCMux32_inw1),
.DataIn_2(MEMOCMux32_inw2),
.DataIn_3(MEMOCMux32_inw3),
.DataIn_4(MEMOCMux32_inw4),
.DataIn_5(MEMOCMux32_inw5),
.DataIn_6(MEMOCMux32_inw6),
.DataIn_7(MEMOCMux32_inw7),
.DataIn_8(MEMOCMux32_inw8),
.DataIn_9(MEMOCMux32_inw9),
.DataIn_10(MEMOCMux32_inw10),
.DataOut_1(MEMOCMux32_outw1),
.sel(MEMOCMux32_selw));
defparam MEMOCMux32.Mux_BW = 32;
assign MEMC32_data_from_Core = MEMOCMux32_outw1;
assign MEMOCMux32_inw1 = dataOutW[31:0]; 
assign MEMOCMux32_inw2 = dataOutW[63:32]; 
assign MEMOCMux32_inw3 = dataOutW[95:64]; 
assign MEMOCMux32_inw4 = dataOutW[127:96]; 
assign MEMOCMux32_inw5 = dataOutW[159:128]; 
assign MEMOCMux32_inw6 = dataOutW[191:160]; 
assign MEMOCMux32_inw7 = dataOutW[223:192]; 
assign MEMOCMux32_inw8 = dataOutW[255:224]; 
assign MEMOCMux32_inw9 = dataOutW[287:256]; 
assign MEMOCMux32_inw10 = globalDataIn[1055:1024]; 
assign MEMOCMux32_selw = mOutConfigW[131:128]; 
assign MEMC32_data_out_ctx2 = mDataFromMem[1055:1024]; 
assign mDataToMem[1055:1024] = MEMC32_data_in_ctx1; 
assign globalDataOut[1055:1024] = MEMC32_data_to_Core; 
assign MEMC32_valid_ctx1 = valid1[32:32]; 
assign MEMC32_write_en_ctx1 = WEn1[32:32]; 
assign MEMC32_stride_ctx1 = stride1[32:32]; 
assign MEMC32_start_addr_ctx1 = startAddr1[197:192]; 
assign MEMC32_burst_count_ctx1 = count1[230:224]; 
assign mAddr1[197:192] = MEMC32_addr_out_ctx1; 
assign mEn1[32:32] = MEMC32_mem_en_ctx1; 
assign mWEn1[32:32] = MEMC32_write_mem_en_ctx1; 
assign MEMC32_valid_ctx2 = valid2[32:32]; 
assign MEMC32_write_en_ctx2 = WEn2[32:32]; 
assign MEMC32_stride_ctx2 = stride2[32:32]; 
assign MEMC32_start_addr_ctx2 = startAddr2[197:192]; 
assign mAddr2[197:192] = MEMC32_addr_out_ctx2; 
assign MEMC32_burst_count_ctx2 = count2[230:224]; 
assign mEn2[32:32] = MEMC32_mem_en_ctx2; 
assign mWEn2[32:32] = MEMC32_write_mem_en_ctx2; 
wire [31:0] MEMOCMux33_inw1;
wire [31:0] MEMOCMux33_inw2;
wire [31:0] MEMOCMux33_inw3;
wire [31:0] MEMOCMux33_inw4;
wire [31:0] MEMOCMux33_inw5;
wire [31:0] MEMOCMux33_inw6;
wire [31:0] MEMOCMux33_inw7;
wire [31:0] MEMOCMux33_inw8;
wire [31:0] MEMOCMux33_inw9;
wire [31:0] MEMOCMux33_inw10;
wire [31:0] MEMOCMux33_outw1;
wire [3:0] MEMOCMux33_selw;
HA_10IM MEMOCMux33 (
.DataIn_1(MEMOCMux33_inw1),
.DataIn_2(MEMOCMux33_inw2),
.DataIn_3(MEMOCMux33_inw3),
.DataIn_4(MEMOCMux33_inw4),
.DataIn_5(MEMOCMux33_inw5),
.DataIn_6(MEMOCMux33_inw6),
.DataIn_7(MEMOCMux33_inw7),
.DataIn_8(MEMOCMux33_inw8),
.DataIn_9(MEMOCMux33_inw9),
.DataIn_10(MEMOCMux33_inw10),
.DataOut_1(MEMOCMux33_outw1),
.sel(MEMOCMux33_selw));
defparam MEMOCMux33.Mux_BW = 32;
assign MEMC33_data_from_Core = MEMOCMux33_outw1;
assign MEMOCMux33_inw1 = dataOutW[31:0]; 
assign MEMOCMux33_inw2 = dataOutW[63:32]; 
assign MEMOCMux33_inw3 = dataOutW[95:64]; 
assign MEMOCMux33_inw4 = dataOutW[127:96]; 
assign MEMOCMux33_inw5 = dataOutW[159:128]; 
assign MEMOCMux33_inw6 = dataOutW[191:160]; 
assign MEMOCMux33_inw7 = dataOutW[223:192]; 
assign MEMOCMux33_inw8 = dataOutW[255:224]; 
assign MEMOCMux33_inw9 = dataOutW[287:256]; 
assign MEMOCMux33_inw10 = globalDataIn[1087:1056]; 
assign MEMOCMux33_selw = mOutConfigW[135:132]; 
assign MEMC33_data_out_ctx2 = mDataFromMem[1087:1056]; 
assign mDataToMem[1087:1056] = MEMC33_data_in_ctx1; 
assign globalDataOut[1087:1056] = MEMC33_data_to_Core; 
assign MEMC33_valid_ctx1 = valid1[33:33]; 
assign MEMC33_write_en_ctx1 = WEn1[33:33]; 
assign MEMC33_stride_ctx1 = stride1[33:33]; 
assign MEMC33_start_addr_ctx1 = startAddr1[203:198]; 
assign MEMC33_burst_count_ctx1 = count1[237:231]; 
assign mAddr1[203:198] = MEMC33_addr_out_ctx1; 
assign mEn1[33:33] = MEMC33_mem_en_ctx1; 
assign mWEn1[33:33] = MEMC33_write_mem_en_ctx1; 
assign MEMC33_valid_ctx2 = valid2[33:33]; 
assign MEMC33_write_en_ctx2 = WEn2[33:33]; 
assign MEMC33_stride_ctx2 = stride2[33:33]; 
assign MEMC33_start_addr_ctx2 = startAddr2[203:198]; 
assign mAddr2[203:198] = MEMC33_addr_out_ctx2; 
assign MEMC33_burst_count_ctx2 = count2[237:231]; 
assign mEn2[33:33] = MEMC33_mem_en_ctx2; 
assign mWEn2[33:33] = MEMC33_write_mem_en_ctx2; 
wire [31:0] MEMOCMux34_inw1;
wire [31:0] MEMOCMux34_inw2;
wire [31:0] MEMOCMux34_inw3;
wire [31:0] MEMOCMux34_inw4;
wire [31:0] MEMOCMux34_inw5;
wire [31:0] MEMOCMux34_inw6;
wire [31:0] MEMOCMux34_inw7;
wire [31:0] MEMOCMux34_inw8;
wire [31:0] MEMOCMux34_inw9;
wire [31:0] MEMOCMux34_inw10;
wire [31:0] MEMOCMux34_outw1;
wire [3:0] MEMOCMux34_selw;
HA_10IM MEMOCMux34 (
.DataIn_1(MEMOCMux34_inw1),
.DataIn_2(MEMOCMux34_inw2),
.DataIn_3(MEMOCMux34_inw3),
.DataIn_4(MEMOCMux34_inw4),
.DataIn_5(MEMOCMux34_inw5),
.DataIn_6(MEMOCMux34_inw6),
.DataIn_7(MEMOCMux34_inw7),
.DataIn_8(MEMOCMux34_inw8),
.DataIn_9(MEMOCMux34_inw9),
.DataIn_10(MEMOCMux34_inw10),
.DataOut_1(MEMOCMux34_outw1),
.sel(MEMOCMux34_selw));
defparam MEMOCMux34.Mux_BW = 32;
assign MEMC34_data_from_Core = MEMOCMux34_outw1;
assign MEMOCMux34_inw1 = dataOutW[31:0]; 
assign MEMOCMux34_inw2 = dataOutW[63:32]; 
assign MEMOCMux34_inw3 = dataOutW[95:64]; 
assign MEMOCMux34_inw4 = dataOutW[127:96]; 
assign MEMOCMux34_inw5 = dataOutW[159:128]; 
assign MEMOCMux34_inw6 = dataOutW[191:160]; 
assign MEMOCMux34_inw7 = dataOutW[223:192]; 
assign MEMOCMux34_inw8 = dataOutW[255:224]; 
assign MEMOCMux34_inw9 = dataOutW[287:256]; 
assign MEMOCMux34_inw10 = globalDataIn[1119:1088]; 
assign MEMOCMux34_selw = mOutConfigW[139:136]; 
assign MEMC34_data_out_ctx2 = mDataFromMem[1119:1088]; 
assign mDataToMem[1119:1088] = MEMC34_data_in_ctx1; 
assign globalDataOut[1119:1088] = MEMC34_data_to_Core; 
assign MEMC34_valid_ctx1 = valid1[34:34]; 
assign MEMC34_write_en_ctx1 = WEn1[34:34]; 
assign MEMC34_stride_ctx1 = stride1[34:34]; 
assign MEMC34_start_addr_ctx1 = startAddr1[209:204]; 
assign MEMC34_burst_count_ctx1 = count1[244:238]; 
assign mAddr1[209:204] = MEMC34_addr_out_ctx1; 
assign mEn1[34:34] = MEMC34_mem_en_ctx1; 
assign mWEn1[34:34] = MEMC34_write_mem_en_ctx1; 
assign MEMC34_valid_ctx2 = valid2[34:34]; 
assign MEMC34_write_en_ctx2 = WEn2[34:34]; 
assign MEMC34_stride_ctx2 = stride2[34:34]; 
assign MEMC34_start_addr_ctx2 = startAddr2[209:204]; 
assign mAddr2[209:204] = MEMC34_addr_out_ctx2; 
assign MEMC34_burst_count_ctx2 = count2[244:238]; 
assign mEn2[34:34] = MEMC34_mem_en_ctx2; 
assign mWEn2[34:34] = MEMC34_write_mem_en_ctx2; 
wire [31:0] MEMOCMux35_inw1;
wire [31:0] MEMOCMux35_inw2;
wire [31:0] MEMOCMux35_inw3;
wire [31:0] MEMOCMux35_inw4;
wire [31:0] MEMOCMux35_inw5;
wire [31:0] MEMOCMux35_inw6;
wire [31:0] MEMOCMux35_inw7;
wire [31:0] MEMOCMux35_inw8;
wire [31:0] MEMOCMux35_inw9;
wire [31:0] MEMOCMux35_inw10;
wire [31:0] MEMOCMux35_outw1;
wire [3:0] MEMOCMux35_selw;
HA_10IM MEMOCMux35 (
.DataIn_1(MEMOCMux35_inw1),
.DataIn_2(MEMOCMux35_inw2),
.DataIn_3(MEMOCMux35_inw3),
.DataIn_4(MEMOCMux35_inw4),
.DataIn_5(MEMOCMux35_inw5),
.DataIn_6(MEMOCMux35_inw6),
.DataIn_7(MEMOCMux35_inw7),
.DataIn_8(MEMOCMux35_inw8),
.DataIn_9(MEMOCMux35_inw9),
.DataIn_10(MEMOCMux35_inw10),
.DataOut_1(MEMOCMux35_outw1),
.sel(MEMOCMux35_selw));
defparam MEMOCMux35.Mux_BW = 32;
assign MEMC35_data_from_Core = MEMOCMux35_outw1;
assign MEMOCMux35_inw1 = dataOutW[31:0]; 
assign MEMOCMux35_inw2 = dataOutW[63:32]; 
assign MEMOCMux35_inw3 = dataOutW[95:64]; 
assign MEMOCMux35_inw4 = dataOutW[127:96]; 
assign MEMOCMux35_inw5 = dataOutW[159:128]; 
assign MEMOCMux35_inw6 = dataOutW[191:160]; 
assign MEMOCMux35_inw7 = dataOutW[223:192]; 
assign MEMOCMux35_inw8 = dataOutW[255:224]; 
assign MEMOCMux35_inw9 = dataOutW[287:256]; 
assign MEMOCMux35_inw10 = globalDataIn[1151:1120]; 
assign MEMOCMux35_selw = mOutConfigW[143:140]; 
assign MEMC35_data_out_ctx2 = mDataFromMem[1151:1120]; 
assign mDataToMem[1151:1120] = MEMC35_data_in_ctx1; 
assign globalDataOut[1151:1120] = MEMC35_data_to_Core; 
assign MEMC35_valid_ctx1 = valid1[35:35]; 
assign MEMC35_write_en_ctx1 = WEn1[35:35]; 
assign MEMC35_stride_ctx1 = stride1[35:35]; 
assign MEMC35_start_addr_ctx1 = startAddr1[215:210]; 
assign MEMC35_burst_count_ctx1 = count1[251:245]; 
assign mAddr1[215:210] = MEMC35_addr_out_ctx1; 
assign mEn1[35:35] = MEMC35_mem_en_ctx1; 
assign mWEn1[35:35] = MEMC35_write_mem_en_ctx1; 
assign MEMC35_valid_ctx2 = valid2[35:35]; 
assign MEMC35_write_en_ctx2 = WEn2[35:35]; 
assign MEMC35_stride_ctx2 = stride2[35:35]; 
assign MEMC35_start_addr_ctx2 = startAddr2[215:210]; 
assign mAddr2[215:210] = MEMC35_addr_out_ctx2; 
assign MEMC35_burst_count_ctx2 = count2[251:245]; 
assign mEn2[35:35] = MEMC35_mem_en_ctx2; 
assign mWEn2[35:35] = MEMC35_write_mem_en_ctx2; 
wire [31:0] MEMOCMux36_inw1;
wire [31:0] MEMOCMux36_inw2;
wire [31:0] MEMOCMux36_inw3;
wire [31:0] MEMOCMux36_inw4;
wire [31:0] MEMOCMux36_inw5;
wire [31:0] MEMOCMux36_inw6;
wire [31:0] MEMOCMux36_inw7;
wire [31:0] MEMOCMux36_inw8;
wire [31:0] MEMOCMux36_inw9;
wire [31:0] MEMOCMux36_inw10;
wire [31:0] MEMOCMux36_outw1;
wire [3:0] MEMOCMux36_selw;
HA_10IM MEMOCMux36 (
.DataIn_1(MEMOCMux36_inw1),
.DataIn_2(MEMOCMux36_inw2),
.DataIn_3(MEMOCMux36_inw3),
.DataIn_4(MEMOCMux36_inw4),
.DataIn_5(MEMOCMux36_inw5),
.DataIn_6(MEMOCMux36_inw6),
.DataIn_7(MEMOCMux36_inw7),
.DataIn_8(MEMOCMux36_inw8),
.DataIn_9(MEMOCMux36_inw9),
.DataIn_10(MEMOCMux36_inw10),
.DataOut_1(MEMOCMux36_outw1),
.sel(MEMOCMux36_selw));
defparam MEMOCMux36.Mux_BW = 32;
assign MEMC36_data_from_Core = MEMOCMux36_outw1;
assign MEMOCMux36_inw1 = dataOutW[31:0]; 
assign MEMOCMux36_inw2 = dataOutW[63:32]; 
assign MEMOCMux36_inw3 = dataOutW[95:64]; 
assign MEMOCMux36_inw4 = dataOutW[127:96]; 
assign MEMOCMux36_inw5 = dataOutW[159:128]; 
assign MEMOCMux36_inw6 = dataOutW[191:160]; 
assign MEMOCMux36_inw7 = dataOutW[223:192]; 
assign MEMOCMux36_inw8 = dataOutW[255:224]; 
assign MEMOCMux36_inw9 = dataOutW[287:256]; 
assign MEMOCMux36_inw10 = globalDataIn[1183:1152]; 
assign MEMOCMux36_selw = mOutConfigW[147:144]; 
assign MEMC36_data_out_ctx2 = mDataFromMem[1183:1152]; 
assign mDataToMem[1183:1152] = MEMC36_data_in_ctx1; 
assign globalDataOut[1183:1152] = MEMC36_data_to_Core; 
assign MEMC36_valid_ctx1 = valid1[36:36]; 
assign MEMC36_write_en_ctx1 = WEn1[36:36]; 
assign MEMC36_stride_ctx1 = stride1[36:36]; 
assign MEMC36_start_addr_ctx1 = startAddr1[221:216]; 
assign MEMC36_burst_count_ctx1 = count1[258:252]; 
assign mAddr1[221:216] = MEMC36_addr_out_ctx1; 
assign mEn1[36:36] = MEMC36_mem_en_ctx1; 
assign mWEn1[36:36] = MEMC36_write_mem_en_ctx1; 
assign MEMC36_valid_ctx2 = valid2[36:36]; 
assign MEMC36_write_en_ctx2 = WEn2[36:36]; 
assign MEMC36_stride_ctx2 = stride2[36:36]; 
assign MEMC36_start_addr_ctx2 = startAddr2[221:216]; 
assign mAddr2[221:216] = MEMC36_addr_out_ctx2; 
assign MEMC36_burst_count_ctx2 = count2[258:252]; 
assign mEn2[36:36] = MEMC36_mem_en_ctx2; 
assign mWEn2[36:36] = MEMC36_write_mem_en_ctx2; 
wire [31:0] MEMOCMux37_inw1;
wire [31:0] MEMOCMux37_inw2;
wire [31:0] MEMOCMux37_inw3;
wire [31:0] MEMOCMux37_inw4;
wire [31:0] MEMOCMux37_inw5;
wire [31:0] MEMOCMux37_inw6;
wire [31:0] MEMOCMux37_inw7;
wire [31:0] MEMOCMux37_inw8;
wire [31:0] MEMOCMux37_inw9;
wire [31:0] MEMOCMux37_inw10;
wire [31:0] MEMOCMux37_outw1;
wire [3:0] MEMOCMux37_selw;
HA_10IM MEMOCMux37 (
.DataIn_1(MEMOCMux37_inw1),
.DataIn_2(MEMOCMux37_inw2),
.DataIn_3(MEMOCMux37_inw3),
.DataIn_4(MEMOCMux37_inw4),
.DataIn_5(MEMOCMux37_inw5),
.DataIn_6(MEMOCMux37_inw6),
.DataIn_7(MEMOCMux37_inw7),
.DataIn_8(MEMOCMux37_inw8),
.DataIn_9(MEMOCMux37_inw9),
.DataIn_10(MEMOCMux37_inw10),
.DataOut_1(MEMOCMux37_outw1),
.sel(MEMOCMux37_selw));
defparam MEMOCMux37.Mux_BW = 32;
assign MEMC37_data_from_Core = MEMOCMux37_outw1;
assign MEMOCMux37_inw1 = dataOutW[31:0]; 
assign MEMOCMux37_inw2 = dataOutW[63:32]; 
assign MEMOCMux37_inw3 = dataOutW[95:64]; 
assign MEMOCMux37_inw4 = dataOutW[127:96]; 
assign MEMOCMux37_inw5 = dataOutW[159:128]; 
assign MEMOCMux37_inw6 = dataOutW[191:160]; 
assign MEMOCMux37_inw7 = dataOutW[223:192]; 
assign MEMOCMux37_inw8 = dataOutW[255:224]; 
assign MEMOCMux37_inw9 = dataOutW[287:256]; 
assign MEMOCMux37_inw10 = globalDataIn[1215:1184]; 
assign MEMOCMux37_selw = mOutConfigW[151:148]; 
assign MEMC37_data_out_ctx2 = mDataFromMem[1215:1184]; 
assign mDataToMem[1215:1184] = MEMC37_data_in_ctx1; 
assign globalDataOut[1215:1184] = MEMC37_data_to_Core; 
assign MEMC37_valid_ctx1 = valid1[37:37]; 
assign MEMC37_write_en_ctx1 = WEn1[37:37]; 
assign MEMC37_stride_ctx1 = stride1[37:37]; 
assign MEMC37_start_addr_ctx1 = startAddr1[227:222]; 
assign MEMC37_burst_count_ctx1 = count1[265:259]; 
assign mAddr1[227:222] = MEMC37_addr_out_ctx1; 
assign mEn1[37:37] = MEMC37_mem_en_ctx1; 
assign mWEn1[37:37] = MEMC37_write_mem_en_ctx1; 
assign MEMC37_valid_ctx2 = valid2[37:37]; 
assign MEMC37_write_en_ctx2 = WEn2[37:37]; 
assign MEMC37_stride_ctx2 = stride2[37:37]; 
assign MEMC37_start_addr_ctx2 = startAddr2[227:222]; 
assign mAddr2[227:222] = MEMC37_addr_out_ctx2; 
assign MEMC37_burst_count_ctx2 = count2[265:259]; 
assign mEn2[37:37] = MEMC37_mem_en_ctx2; 
assign mWEn2[37:37] = MEMC37_write_mem_en_ctx2; 
wire [31:0] MEMOCMux38_inw1;
wire [31:0] MEMOCMux38_inw2;
wire [31:0] MEMOCMux38_inw3;
wire [31:0] MEMOCMux38_inw4;
wire [31:0] MEMOCMux38_inw5;
wire [31:0] MEMOCMux38_inw6;
wire [31:0] MEMOCMux38_inw7;
wire [31:0] MEMOCMux38_inw8;
wire [31:0] MEMOCMux38_inw9;
wire [31:0] MEMOCMux38_inw10;
wire [31:0] MEMOCMux38_outw1;
wire [3:0] MEMOCMux38_selw;
HA_10IM MEMOCMux38 (
.DataIn_1(MEMOCMux38_inw1),
.DataIn_2(MEMOCMux38_inw2),
.DataIn_3(MEMOCMux38_inw3),
.DataIn_4(MEMOCMux38_inw4),
.DataIn_5(MEMOCMux38_inw5),
.DataIn_6(MEMOCMux38_inw6),
.DataIn_7(MEMOCMux38_inw7),
.DataIn_8(MEMOCMux38_inw8),
.DataIn_9(MEMOCMux38_inw9),
.DataIn_10(MEMOCMux38_inw10),
.DataOut_1(MEMOCMux38_outw1),
.sel(MEMOCMux38_selw));
defparam MEMOCMux38.Mux_BW = 32;
assign MEMC38_data_from_Core = MEMOCMux38_outw1;
assign MEMOCMux38_inw1 = dataOutW[31:0]; 
assign MEMOCMux38_inw2 = dataOutW[63:32]; 
assign MEMOCMux38_inw3 = dataOutW[95:64]; 
assign MEMOCMux38_inw4 = dataOutW[127:96]; 
assign MEMOCMux38_inw5 = dataOutW[159:128]; 
assign MEMOCMux38_inw6 = dataOutW[191:160]; 
assign MEMOCMux38_inw7 = dataOutW[223:192]; 
assign MEMOCMux38_inw8 = dataOutW[255:224]; 
assign MEMOCMux38_inw9 = dataOutW[287:256]; 
assign MEMOCMux38_inw10 = globalDataIn[1247:1216]; 
assign MEMOCMux38_selw = mOutConfigW[155:152]; 
assign MEMC38_data_out_ctx2 = mDataFromMem[1247:1216]; 
assign mDataToMem[1247:1216] = MEMC38_data_in_ctx1; 
assign globalDataOut[1247:1216] = MEMC38_data_to_Core; 
assign MEMC38_valid_ctx1 = valid1[38:38]; 
assign MEMC38_write_en_ctx1 = WEn1[38:38]; 
assign MEMC38_stride_ctx1 = stride1[38:38]; 
assign MEMC38_start_addr_ctx1 = startAddr1[233:228]; 
assign MEMC38_burst_count_ctx1 = count1[272:266]; 
assign mAddr1[233:228] = MEMC38_addr_out_ctx1; 
assign mEn1[38:38] = MEMC38_mem_en_ctx1; 
assign mWEn1[38:38] = MEMC38_write_mem_en_ctx1; 
assign MEMC38_valid_ctx2 = valid2[38:38]; 
assign MEMC38_write_en_ctx2 = WEn2[38:38]; 
assign MEMC38_stride_ctx2 = stride2[38:38]; 
assign MEMC38_start_addr_ctx2 = startAddr2[233:228]; 
assign mAddr2[233:228] = MEMC38_addr_out_ctx2; 
assign MEMC38_burst_count_ctx2 = count2[272:266]; 
assign mEn2[38:38] = MEMC38_mem_en_ctx2; 
assign mWEn2[38:38] = MEMC38_write_mem_en_ctx2; 
wire [31:0] MEMOCMux39_inw1;
wire [31:0] MEMOCMux39_inw2;
wire [31:0] MEMOCMux39_inw3;
wire [31:0] MEMOCMux39_inw4;
wire [31:0] MEMOCMux39_inw5;
wire [31:0] MEMOCMux39_inw6;
wire [31:0] MEMOCMux39_inw7;
wire [31:0] MEMOCMux39_inw8;
wire [31:0] MEMOCMux39_inw9;
wire [31:0] MEMOCMux39_inw10;
wire [31:0] MEMOCMux39_outw1;
wire [3:0] MEMOCMux39_selw;
HA_10IM MEMOCMux39 (
.DataIn_1(MEMOCMux39_inw1),
.DataIn_2(MEMOCMux39_inw2),
.DataIn_3(MEMOCMux39_inw3),
.DataIn_4(MEMOCMux39_inw4),
.DataIn_5(MEMOCMux39_inw5),
.DataIn_6(MEMOCMux39_inw6),
.DataIn_7(MEMOCMux39_inw7),
.DataIn_8(MEMOCMux39_inw8),
.DataIn_9(MEMOCMux39_inw9),
.DataIn_10(MEMOCMux39_inw10),
.DataOut_1(MEMOCMux39_outw1),
.sel(MEMOCMux39_selw));
defparam MEMOCMux39.Mux_BW = 32;
assign MEMC39_data_from_Core = MEMOCMux39_outw1;
assign MEMOCMux39_inw1 = dataOutW[31:0]; 
assign MEMOCMux39_inw2 = dataOutW[63:32]; 
assign MEMOCMux39_inw3 = dataOutW[95:64]; 
assign MEMOCMux39_inw4 = dataOutW[127:96]; 
assign MEMOCMux39_inw5 = dataOutW[159:128]; 
assign MEMOCMux39_inw6 = dataOutW[191:160]; 
assign MEMOCMux39_inw7 = dataOutW[223:192]; 
assign MEMOCMux39_inw8 = dataOutW[255:224]; 
assign MEMOCMux39_inw9 = dataOutW[287:256]; 
assign MEMOCMux39_inw10 = globalDataIn[1279:1248]; 
assign MEMOCMux39_selw = mOutConfigW[159:156]; 
assign MEMC39_data_out_ctx2 = mDataFromMem[1279:1248]; 
assign mDataToMem[1279:1248] = MEMC39_data_in_ctx1; 
assign globalDataOut[1279:1248] = MEMC39_data_to_Core; 
assign MEMC39_valid_ctx1 = valid1[39:39]; 
assign MEMC39_write_en_ctx1 = WEn1[39:39]; 
assign MEMC39_stride_ctx1 = stride1[39:39]; 
assign MEMC39_start_addr_ctx1 = startAddr1[239:234]; 
assign MEMC39_burst_count_ctx1 = count1[279:273]; 
assign mAddr1[239:234] = MEMC39_addr_out_ctx1; 
assign mEn1[39:39] = MEMC39_mem_en_ctx1; 
assign mWEn1[39:39] = MEMC39_write_mem_en_ctx1; 
assign MEMC39_valid_ctx2 = valid2[39:39]; 
assign MEMC39_write_en_ctx2 = WEn2[39:39]; 
assign MEMC39_stride_ctx2 = stride2[39:39]; 
assign MEMC39_start_addr_ctx2 = startAddr2[239:234]; 
assign mAddr2[239:234] = MEMC39_addr_out_ctx2; 
assign MEMC39_burst_count_ctx2 = count2[279:273]; 
assign mEn2[39:39] = MEMC39_mem_en_ctx2; 
assign mWEn2[39:39] = MEMC39_write_mem_en_ctx2; 
wire [31:0] MEMOCMux40_inw1;
wire [31:0] MEMOCMux40_inw2;
wire [31:0] MEMOCMux40_inw3;
wire [31:0] MEMOCMux40_inw4;
wire [31:0] MEMOCMux40_inw5;
wire [31:0] MEMOCMux40_inw6;
wire [31:0] MEMOCMux40_inw7;
wire [31:0] MEMOCMux40_inw8;
wire [31:0] MEMOCMux40_inw9;
wire [31:0] MEMOCMux40_inw10;
wire [31:0] MEMOCMux40_outw1;
wire [3:0] MEMOCMux40_selw;
HA_10IM MEMOCMux40 (
.DataIn_1(MEMOCMux40_inw1),
.DataIn_2(MEMOCMux40_inw2),
.DataIn_3(MEMOCMux40_inw3),
.DataIn_4(MEMOCMux40_inw4),
.DataIn_5(MEMOCMux40_inw5),
.DataIn_6(MEMOCMux40_inw6),
.DataIn_7(MEMOCMux40_inw7),
.DataIn_8(MEMOCMux40_inw8),
.DataIn_9(MEMOCMux40_inw9),
.DataIn_10(MEMOCMux40_inw10),
.DataOut_1(MEMOCMux40_outw1),
.sel(MEMOCMux40_selw));
defparam MEMOCMux40.Mux_BW = 32;
assign MEMC40_data_from_Core = MEMOCMux40_outw1;
assign MEMOCMux40_inw1 = dataOutW[31:0]; 
assign MEMOCMux40_inw2 = dataOutW[63:32]; 
assign MEMOCMux40_inw3 = dataOutW[95:64]; 
assign MEMOCMux40_inw4 = dataOutW[127:96]; 
assign MEMOCMux40_inw5 = dataOutW[159:128]; 
assign MEMOCMux40_inw6 = dataOutW[191:160]; 
assign MEMOCMux40_inw7 = dataOutW[223:192]; 
assign MEMOCMux40_inw8 = dataOutW[255:224]; 
assign MEMOCMux40_inw9 = dataOutW[287:256]; 
assign MEMOCMux40_inw10 = globalDataIn[1311:1280]; 
assign MEMOCMux40_selw = mOutConfigW[163:160]; 
assign MEMC40_data_out_ctx2 = mDataFromMem[1311:1280]; 
assign mDataToMem[1311:1280] = MEMC40_data_in_ctx1; 
assign globalDataOut[1311:1280] = MEMC40_data_to_Core; 
assign MEMC40_valid_ctx1 = valid1[40:40]; 
assign MEMC40_write_en_ctx1 = WEn1[40:40]; 
assign MEMC40_stride_ctx1 = stride1[40:40]; 
assign MEMC40_start_addr_ctx1 = startAddr1[245:240]; 
assign MEMC40_burst_count_ctx1 = count1[286:280]; 
assign mAddr1[245:240] = MEMC40_addr_out_ctx1; 
assign mEn1[40:40] = MEMC40_mem_en_ctx1; 
assign mWEn1[40:40] = MEMC40_write_mem_en_ctx1; 
assign MEMC40_valid_ctx2 = valid2[40:40]; 
assign MEMC40_write_en_ctx2 = WEn2[40:40]; 
assign MEMC40_stride_ctx2 = stride2[40:40]; 
assign MEMC40_start_addr_ctx2 = startAddr2[245:240]; 
assign mAddr2[245:240] = MEMC40_addr_out_ctx2; 
assign MEMC40_burst_count_ctx2 = count2[286:280]; 
assign mEn2[40:40] = MEMC40_mem_en_ctx2; 
assign mWEn2[40:40] = MEMC40_write_mem_en_ctx2; 
wire [31:0] MEMOCMux41_inw1;
wire [31:0] MEMOCMux41_inw2;
wire [31:0] MEMOCMux41_inw3;
wire [31:0] MEMOCMux41_inw4;
wire [31:0] MEMOCMux41_inw5;
wire [31:0] MEMOCMux41_inw6;
wire [31:0] MEMOCMux41_inw7;
wire [31:0] MEMOCMux41_inw8;
wire [31:0] MEMOCMux41_inw9;
wire [31:0] MEMOCMux41_inw10;
wire [31:0] MEMOCMux41_outw1;
wire [3:0] MEMOCMux41_selw;
HA_10IM MEMOCMux41 (
.DataIn_1(MEMOCMux41_inw1),
.DataIn_2(MEMOCMux41_inw2),
.DataIn_3(MEMOCMux41_inw3),
.DataIn_4(MEMOCMux41_inw4),
.DataIn_5(MEMOCMux41_inw5),
.DataIn_6(MEMOCMux41_inw6),
.DataIn_7(MEMOCMux41_inw7),
.DataIn_8(MEMOCMux41_inw8),
.DataIn_9(MEMOCMux41_inw9),
.DataIn_10(MEMOCMux41_inw10),
.DataOut_1(MEMOCMux41_outw1),
.sel(MEMOCMux41_selw));
defparam MEMOCMux41.Mux_BW = 32;
assign MEMC41_data_from_Core = MEMOCMux41_outw1;
assign MEMOCMux41_inw1 = dataOutW[31:0]; 
assign MEMOCMux41_inw2 = dataOutW[63:32]; 
assign MEMOCMux41_inw3 = dataOutW[95:64]; 
assign MEMOCMux41_inw4 = dataOutW[127:96]; 
assign MEMOCMux41_inw5 = dataOutW[159:128]; 
assign MEMOCMux41_inw6 = dataOutW[191:160]; 
assign MEMOCMux41_inw7 = dataOutW[223:192]; 
assign MEMOCMux41_inw8 = dataOutW[255:224]; 
assign MEMOCMux41_inw9 = dataOutW[287:256]; 
assign MEMOCMux41_inw10 = globalDataIn[1343:1312]; 
assign MEMOCMux41_selw = mOutConfigW[167:164]; 
assign MEMC41_data_out_ctx2 = mDataFromMem[1343:1312]; 
assign mDataToMem[1343:1312] = MEMC41_data_in_ctx1; 
assign globalDataOut[1343:1312] = MEMC41_data_to_Core; 
assign MEMC41_valid_ctx1 = valid1[41:41]; 
assign MEMC41_write_en_ctx1 = WEn1[41:41]; 
assign MEMC41_stride_ctx1 = stride1[41:41]; 
assign MEMC41_start_addr_ctx1 = startAddr1[251:246]; 
assign MEMC41_burst_count_ctx1 = count1[293:287]; 
assign mAddr1[251:246] = MEMC41_addr_out_ctx1; 
assign mEn1[41:41] = MEMC41_mem_en_ctx1; 
assign mWEn1[41:41] = MEMC41_write_mem_en_ctx1; 
assign MEMC41_valid_ctx2 = valid2[41:41]; 
assign MEMC41_write_en_ctx2 = WEn2[41:41]; 
assign MEMC41_stride_ctx2 = stride2[41:41]; 
assign MEMC41_start_addr_ctx2 = startAddr2[251:246]; 
assign mAddr2[251:246] = MEMC41_addr_out_ctx2; 
assign MEMC41_burst_count_ctx2 = count2[293:287]; 
assign mEn2[41:41] = MEMC41_mem_en_ctx2; 
assign mWEn2[41:41] = MEMC41_write_mem_en_ctx2; 
wire [31:0] MEMOCMux42_inw1;
wire [31:0] MEMOCMux42_inw2;
wire [31:0] MEMOCMux42_inw3;
wire [31:0] MEMOCMux42_inw4;
wire [31:0] MEMOCMux42_inw5;
wire [31:0] MEMOCMux42_inw6;
wire [31:0] MEMOCMux42_inw7;
wire [31:0] MEMOCMux42_inw8;
wire [31:0] MEMOCMux42_inw9;
wire [31:0] MEMOCMux42_inw10;
wire [31:0] MEMOCMux42_outw1;
wire [3:0] MEMOCMux42_selw;
HA_10IM MEMOCMux42 (
.DataIn_1(MEMOCMux42_inw1),
.DataIn_2(MEMOCMux42_inw2),
.DataIn_3(MEMOCMux42_inw3),
.DataIn_4(MEMOCMux42_inw4),
.DataIn_5(MEMOCMux42_inw5),
.DataIn_6(MEMOCMux42_inw6),
.DataIn_7(MEMOCMux42_inw7),
.DataIn_8(MEMOCMux42_inw8),
.DataIn_9(MEMOCMux42_inw9),
.DataIn_10(MEMOCMux42_inw10),
.DataOut_1(MEMOCMux42_outw1),
.sel(MEMOCMux42_selw));
defparam MEMOCMux42.Mux_BW = 32;
assign MEMC42_data_from_Core = MEMOCMux42_outw1;
assign MEMOCMux42_inw1 = dataOutW[31:0]; 
assign MEMOCMux42_inw2 = dataOutW[63:32]; 
assign MEMOCMux42_inw3 = dataOutW[95:64]; 
assign MEMOCMux42_inw4 = dataOutW[127:96]; 
assign MEMOCMux42_inw5 = dataOutW[159:128]; 
assign MEMOCMux42_inw6 = dataOutW[191:160]; 
assign MEMOCMux42_inw7 = dataOutW[223:192]; 
assign MEMOCMux42_inw8 = dataOutW[255:224]; 
assign MEMOCMux42_inw9 = dataOutW[287:256]; 
assign MEMOCMux42_inw10 = globalDataIn[1375:1344]; 
assign MEMOCMux42_selw = mOutConfigW[171:168]; 
assign MEMC42_data_out_ctx2 = mDataFromMem[1375:1344]; 
assign mDataToMem[1375:1344] = MEMC42_data_in_ctx1; 
assign globalDataOut[1375:1344] = MEMC42_data_to_Core; 
assign MEMC42_valid_ctx1 = valid1[42:42]; 
assign MEMC42_write_en_ctx1 = WEn1[42:42]; 
assign MEMC42_stride_ctx1 = stride1[42:42]; 
assign MEMC42_start_addr_ctx1 = startAddr1[257:252]; 
assign MEMC42_burst_count_ctx1 = count1[300:294]; 
assign mAddr1[257:252] = MEMC42_addr_out_ctx1; 
assign mEn1[42:42] = MEMC42_mem_en_ctx1; 
assign mWEn1[42:42] = MEMC42_write_mem_en_ctx1; 
assign MEMC42_valid_ctx2 = valid2[42:42]; 
assign MEMC42_write_en_ctx2 = WEn2[42:42]; 
assign MEMC42_stride_ctx2 = stride2[42:42]; 
assign MEMC42_start_addr_ctx2 = startAddr2[257:252]; 
assign mAddr2[257:252] = MEMC42_addr_out_ctx2; 
assign MEMC42_burst_count_ctx2 = count2[300:294]; 
assign mEn2[42:42] = MEMC42_mem_en_ctx2; 
assign mWEn2[42:42] = MEMC42_write_mem_en_ctx2; 
wire [31:0] MEMOCMux43_inw1;
wire [31:0] MEMOCMux43_inw2;
wire [31:0] MEMOCMux43_inw3;
wire [31:0] MEMOCMux43_inw4;
wire [31:0] MEMOCMux43_inw5;
wire [31:0] MEMOCMux43_inw6;
wire [31:0] MEMOCMux43_inw7;
wire [31:0] MEMOCMux43_inw8;
wire [31:0] MEMOCMux43_inw9;
wire [31:0] MEMOCMux43_inw10;
wire [31:0] MEMOCMux43_outw1;
wire [3:0] MEMOCMux43_selw;
HA_10IM MEMOCMux43 (
.DataIn_1(MEMOCMux43_inw1),
.DataIn_2(MEMOCMux43_inw2),
.DataIn_3(MEMOCMux43_inw3),
.DataIn_4(MEMOCMux43_inw4),
.DataIn_5(MEMOCMux43_inw5),
.DataIn_6(MEMOCMux43_inw6),
.DataIn_7(MEMOCMux43_inw7),
.DataIn_8(MEMOCMux43_inw8),
.DataIn_9(MEMOCMux43_inw9),
.DataIn_10(MEMOCMux43_inw10),
.DataOut_1(MEMOCMux43_outw1),
.sel(MEMOCMux43_selw));
defparam MEMOCMux43.Mux_BW = 32;
assign MEMC43_data_from_Core = MEMOCMux43_outw1;
assign MEMOCMux43_inw1 = dataOutW[31:0]; 
assign MEMOCMux43_inw2 = dataOutW[63:32]; 
assign MEMOCMux43_inw3 = dataOutW[95:64]; 
assign MEMOCMux43_inw4 = dataOutW[127:96]; 
assign MEMOCMux43_inw5 = dataOutW[159:128]; 
assign MEMOCMux43_inw6 = dataOutW[191:160]; 
assign MEMOCMux43_inw7 = dataOutW[223:192]; 
assign MEMOCMux43_inw8 = dataOutW[255:224]; 
assign MEMOCMux43_inw9 = dataOutW[287:256]; 
assign MEMOCMux43_inw10 = globalDataIn[1407:1376]; 
assign MEMOCMux43_selw = mOutConfigW[175:172]; 
assign MEMC43_data_out_ctx2 = mDataFromMem[1407:1376]; 
assign mDataToMem[1407:1376] = MEMC43_data_in_ctx1; 
assign globalDataOut[1407:1376] = MEMC43_data_to_Core; 
assign MEMC43_valid_ctx1 = valid1[43:43]; 
assign MEMC43_write_en_ctx1 = WEn1[43:43]; 
assign MEMC43_stride_ctx1 = stride1[43:43]; 
assign MEMC43_start_addr_ctx1 = startAddr1[263:258]; 
assign MEMC43_burst_count_ctx1 = count1[307:301]; 
assign mAddr1[263:258] = MEMC43_addr_out_ctx1; 
assign mEn1[43:43] = MEMC43_mem_en_ctx1; 
assign mWEn1[43:43] = MEMC43_write_mem_en_ctx1; 
assign MEMC43_valid_ctx2 = valid2[43:43]; 
assign MEMC43_write_en_ctx2 = WEn2[43:43]; 
assign MEMC43_stride_ctx2 = stride2[43:43]; 
assign MEMC43_start_addr_ctx2 = startAddr2[263:258]; 
assign mAddr2[263:258] = MEMC43_addr_out_ctx2; 
assign MEMC43_burst_count_ctx2 = count2[307:301]; 
assign mEn2[43:43] = MEMC43_mem_en_ctx2; 
assign mWEn2[43:43] = MEMC43_write_mem_en_ctx2; 
wire [31:0] MEMOCMux44_inw1;
wire [31:0] MEMOCMux44_inw2;
wire [31:0] MEMOCMux44_inw3;
wire [31:0] MEMOCMux44_inw4;
wire [31:0] MEMOCMux44_inw5;
wire [31:0] MEMOCMux44_inw6;
wire [31:0] MEMOCMux44_inw7;
wire [31:0] MEMOCMux44_inw8;
wire [31:0] MEMOCMux44_inw9;
wire [31:0] MEMOCMux44_inw10;
wire [31:0] MEMOCMux44_outw1;
wire [3:0] MEMOCMux44_selw;
HA_10IM MEMOCMux44 (
.DataIn_1(MEMOCMux44_inw1),
.DataIn_2(MEMOCMux44_inw2),
.DataIn_3(MEMOCMux44_inw3),
.DataIn_4(MEMOCMux44_inw4),
.DataIn_5(MEMOCMux44_inw5),
.DataIn_6(MEMOCMux44_inw6),
.DataIn_7(MEMOCMux44_inw7),
.DataIn_8(MEMOCMux44_inw8),
.DataIn_9(MEMOCMux44_inw9),
.DataIn_10(MEMOCMux44_inw10),
.DataOut_1(MEMOCMux44_outw1),
.sel(MEMOCMux44_selw));
defparam MEMOCMux44.Mux_BW = 32;
assign MEMC44_data_from_Core = MEMOCMux44_outw1;
assign MEMOCMux44_inw1 = dataOutW[31:0]; 
assign MEMOCMux44_inw2 = dataOutW[63:32]; 
assign MEMOCMux44_inw3 = dataOutW[95:64]; 
assign MEMOCMux44_inw4 = dataOutW[127:96]; 
assign MEMOCMux44_inw5 = dataOutW[159:128]; 
assign MEMOCMux44_inw6 = dataOutW[191:160]; 
assign MEMOCMux44_inw7 = dataOutW[223:192]; 
assign MEMOCMux44_inw8 = dataOutW[255:224]; 
assign MEMOCMux44_inw9 = dataOutW[287:256]; 
assign MEMOCMux44_inw10 = globalDataIn[1439:1408]; 
assign MEMOCMux44_selw = mOutConfigW[179:176]; 
assign MEMC44_data_out_ctx2 = mDataFromMem[1439:1408]; 
assign mDataToMem[1439:1408] = MEMC44_data_in_ctx1; 
assign globalDataOut[1439:1408] = MEMC44_data_to_Core; 
assign MEMC44_valid_ctx1 = valid1[44:44]; 
assign MEMC44_write_en_ctx1 = WEn1[44:44]; 
assign MEMC44_stride_ctx1 = stride1[44:44]; 
assign MEMC44_start_addr_ctx1 = startAddr1[269:264]; 
assign MEMC44_burst_count_ctx1 = count1[314:308]; 
assign mAddr1[269:264] = MEMC44_addr_out_ctx1; 
assign mEn1[44:44] = MEMC44_mem_en_ctx1; 
assign mWEn1[44:44] = MEMC44_write_mem_en_ctx1; 
assign MEMC44_valid_ctx2 = valid2[44:44]; 
assign MEMC44_write_en_ctx2 = WEn2[44:44]; 
assign MEMC44_stride_ctx2 = stride2[44:44]; 
assign MEMC44_start_addr_ctx2 = startAddr2[269:264]; 
assign mAddr2[269:264] = MEMC44_addr_out_ctx2; 
assign MEMC44_burst_count_ctx2 = count2[314:308]; 
assign mEn2[44:44] = MEMC44_mem_en_ctx2; 
assign mWEn2[44:44] = MEMC44_write_mem_en_ctx2; 
wire [31:0] MEMOCMux45_inw1;
wire [31:0] MEMOCMux45_inw2;
wire [31:0] MEMOCMux45_inw3;
wire [31:0] MEMOCMux45_inw4;
wire [31:0] MEMOCMux45_inw5;
wire [31:0] MEMOCMux45_inw6;
wire [31:0] MEMOCMux45_inw7;
wire [31:0] MEMOCMux45_inw8;
wire [31:0] MEMOCMux45_inw9;
wire [31:0] MEMOCMux45_inw10;
wire [31:0] MEMOCMux45_outw1;
wire [3:0] MEMOCMux45_selw;
HA_10IM MEMOCMux45 (
.DataIn_1(MEMOCMux45_inw1),
.DataIn_2(MEMOCMux45_inw2),
.DataIn_3(MEMOCMux45_inw3),
.DataIn_4(MEMOCMux45_inw4),
.DataIn_5(MEMOCMux45_inw5),
.DataIn_6(MEMOCMux45_inw6),
.DataIn_7(MEMOCMux45_inw7),
.DataIn_8(MEMOCMux45_inw8),
.DataIn_9(MEMOCMux45_inw9),
.DataIn_10(MEMOCMux45_inw10),
.DataOut_1(MEMOCMux45_outw1),
.sel(MEMOCMux45_selw));
defparam MEMOCMux45.Mux_BW = 32;
assign MEMC45_data_from_Core = MEMOCMux45_outw1;
assign MEMOCMux45_inw1 = dataOutW[31:0]; 
assign MEMOCMux45_inw2 = dataOutW[63:32]; 
assign MEMOCMux45_inw3 = dataOutW[95:64]; 
assign MEMOCMux45_inw4 = dataOutW[127:96]; 
assign MEMOCMux45_inw5 = dataOutW[159:128]; 
assign MEMOCMux45_inw6 = dataOutW[191:160]; 
assign MEMOCMux45_inw7 = dataOutW[223:192]; 
assign MEMOCMux45_inw8 = dataOutW[255:224]; 
assign MEMOCMux45_inw9 = dataOutW[287:256]; 
assign MEMOCMux45_inw10 = globalDataIn[1471:1440]; 
assign MEMOCMux45_selw = mOutConfigW[183:180]; 
assign MEMC45_data_out_ctx2 = mDataFromMem[1471:1440]; 
assign mDataToMem[1471:1440] = MEMC45_data_in_ctx1; 
assign globalDataOut[1471:1440] = MEMC45_data_to_Core; 
assign MEMC45_valid_ctx1 = valid1[45:45]; 
assign MEMC45_write_en_ctx1 = WEn1[45:45]; 
assign MEMC45_stride_ctx1 = stride1[45:45]; 
assign MEMC45_start_addr_ctx1 = startAddr1[275:270]; 
assign MEMC45_burst_count_ctx1 = count1[321:315]; 
assign mAddr1[275:270] = MEMC45_addr_out_ctx1; 
assign mEn1[45:45] = MEMC45_mem_en_ctx1; 
assign mWEn1[45:45] = MEMC45_write_mem_en_ctx1; 
assign MEMC45_valid_ctx2 = valid2[45:45]; 
assign MEMC45_write_en_ctx2 = WEn2[45:45]; 
assign MEMC45_stride_ctx2 = stride2[45:45]; 
assign MEMC45_start_addr_ctx2 = startAddr2[275:270]; 
assign mAddr2[275:270] = MEMC45_addr_out_ctx2; 
assign MEMC45_burst_count_ctx2 = count2[321:315]; 
assign mEn2[45:45] = MEMC45_mem_en_ctx2; 
assign mWEn2[45:45] = MEMC45_write_mem_en_ctx2; 
wire [31:0] MEMOCMux46_inw1;
wire [31:0] MEMOCMux46_inw2;
wire [31:0] MEMOCMux46_inw3;
wire [31:0] MEMOCMux46_inw4;
wire [31:0] MEMOCMux46_inw5;
wire [31:0] MEMOCMux46_inw6;
wire [31:0] MEMOCMux46_inw7;
wire [31:0] MEMOCMux46_inw8;
wire [31:0] MEMOCMux46_inw9;
wire [31:0] MEMOCMux46_inw10;
wire [31:0] MEMOCMux46_outw1;
wire [3:0] MEMOCMux46_selw;
HA_10IM MEMOCMux46 (
.DataIn_1(MEMOCMux46_inw1),
.DataIn_2(MEMOCMux46_inw2),
.DataIn_3(MEMOCMux46_inw3),
.DataIn_4(MEMOCMux46_inw4),
.DataIn_5(MEMOCMux46_inw5),
.DataIn_6(MEMOCMux46_inw6),
.DataIn_7(MEMOCMux46_inw7),
.DataIn_8(MEMOCMux46_inw8),
.DataIn_9(MEMOCMux46_inw9),
.DataIn_10(MEMOCMux46_inw10),
.DataOut_1(MEMOCMux46_outw1),
.sel(MEMOCMux46_selw));
defparam MEMOCMux46.Mux_BW = 32;
assign MEMC46_data_from_Core = MEMOCMux46_outw1;
assign MEMOCMux46_inw1 = dataOutW[31:0]; 
assign MEMOCMux46_inw2 = dataOutW[63:32]; 
assign MEMOCMux46_inw3 = dataOutW[95:64]; 
assign MEMOCMux46_inw4 = dataOutW[127:96]; 
assign MEMOCMux46_inw5 = dataOutW[159:128]; 
assign MEMOCMux46_inw6 = dataOutW[191:160]; 
assign MEMOCMux46_inw7 = dataOutW[223:192]; 
assign MEMOCMux46_inw8 = dataOutW[255:224]; 
assign MEMOCMux46_inw9 = dataOutW[287:256]; 
assign MEMOCMux46_inw10 = globalDataIn[1503:1472]; 
assign MEMOCMux46_selw = mOutConfigW[187:184]; 
assign MEMC46_data_out_ctx2 = mDataFromMem[1503:1472]; 
assign mDataToMem[1503:1472] = MEMC46_data_in_ctx1; 
assign globalDataOut[1503:1472] = MEMC46_data_to_Core; 
assign MEMC46_valid_ctx1 = valid1[46:46]; 
assign MEMC46_write_en_ctx1 = WEn1[46:46]; 
assign MEMC46_stride_ctx1 = stride1[46:46]; 
assign MEMC46_start_addr_ctx1 = startAddr1[281:276]; 
assign MEMC46_burst_count_ctx1 = count1[328:322]; 
assign mAddr1[281:276] = MEMC46_addr_out_ctx1; 
assign mEn1[46:46] = MEMC46_mem_en_ctx1; 
assign mWEn1[46:46] = MEMC46_write_mem_en_ctx1; 
assign MEMC46_valid_ctx2 = valid2[46:46]; 
assign MEMC46_write_en_ctx2 = WEn2[46:46]; 
assign MEMC46_stride_ctx2 = stride2[46:46]; 
assign MEMC46_start_addr_ctx2 = startAddr2[281:276]; 
assign mAddr2[281:276] = MEMC46_addr_out_ctx2; 
assign MEMC46_burst_count_ctx2 = count2[328:322]; 
assign mEn2[46:46] = MEMC46_mem_en_ctx2; 
assign mWEn2[46:46] = MEMC46_write_mem_en_ctx2; 
wire [31:0] MEMOCMux47_inw1;
wire [31:0] MEMOCMux47_inw2;
wire [31:0] MEMOCMux47_inw3;
wire [31:0] MEMOCMux47_inw4;
wire [31:0] MEMOCMux47_inw5;
wire [31:0] MEMOCMux47_inw6;
wire [31:0] MEMOCMux47_inw7;
wire [31:0] MEMOCMux47_inw8;
wire [31:0] MEMOCMux47_inw9;
wire [31:0] MEMOCMux47_inw10;
wire [31:0] MEMOCMux47_outw1;
wire [3:0] MEMOCMux47_selw;
HA_10IM MEMOCMux47 (
.DataIn_1(MEMOCMux47_inw1),
.DataIn_2(MEMOCMux47_inw2),
.DataIn_3(MEMOCMux47_inw3),
.DataIn_4(MEMOCMux47_inw4),
.DataIn_5(MEMOCMux47_inw5),
.DataIn_6(MEMOCMux47_inw6),
.DataIn_7(MEMOCMux47_inw7),
.DataIn_8(MEMOCMux47_inw8),
.DataIn_9(MEMOCMux47_inw9),
.DataIn_10(MEMOCMux47_inw10),
.DataOut_1(MEMOCMux47_outw1),
.sel(MEMOCMux47_selw));
defparam MEMOCMux47.Mux_BW = 32;
assign MEMC47_data_from_Core = MEMOCMux47_outw1;
assign MEMOCMux47_inw1 = dataOutW[31:0]; 
assign MEMOCMux47_inw2 = dataOutW[63:32]; 
assign MEMOCMux47_inw3 = dataOutW[95:64]; 
assign MEMOCMux47_inw4 = dataOutW[127:96]; 
assign MEMOCMux47_inw5 = dataOutW[159:128]; 
assign MEMOCMux47_inw6 = dataOutW[191:160]; 
assign MEMOCMux47_inw7 = dataOutW[223:192]; 
assign MEMOCMux47_inw8 = dataOutW[255:224]; 
assign MEMOCMux47_inw9 = dataOutW[287:256]; 
assign MEMOCMux47_inw10 = globalDataIn[1535:1504]; 
assign MEMOCMux47_selw = mOutConfigW[191:188]; 
assign MEMC47_data_out_ctx2 = mDataFromMem[1535:1504]; 
assign mDataToMem[1535:1504] = MEMC47_data_in_ctx1; 
assign globalDataOut[1535:1504] = MEMC47_data_to_Core; 
assign MEMC47_valid_ctx1 = valid1[47:47]; 
assign MEMC47_write_en_ctx1 = WEn1[47:47]; 
assign MEMC47_stride_ctx1 = stride1[47:47]; 
assign MEMC47_start_addr_ctx1 = startAddr1[287:282]; 
assign MEMC47_burst_count_ctx1 = count1[335:329]; 
assign mAddr1[287:282] = MEMC47_addr_out_ctx1; 
assign mEn1[47:47] = MEMC47_mem_en_ctx1; 
assign mWEn1[47:47] = MEMC47_write_mem_en_ctx1; 
assign MEMC47_valid_ctx2 = valid2[47:47]; 
assign MEMC47_write_en_ctx2 = WEn2[47:47]; 
assign MEMC47_stride_ctx2 = stride2[47:47]; 
assign MEMC47_start_addr_ctx2 = startAddr2[287:282]; 
assign mAddr2[287:282] = MEMC47_addr_out_ctx2; 
assign MEMC47_burst_count_ctx2 = count2[335:329]; 
assign mEn2[47:47] = MEMC47_mem_en_ctx2; 
assign mWEn2[47:47] = MEMC47_write_mem_en_ctx2; 
wire [31:0] MEMOCMux48_inw1;
wire [31:0] MEMOCMux48_inw2;
wire [31:0] MEMOCMux48_inw3;
wire [31:0] MEMOCMux48_inw4;
wire [31:0] MEMOCMux48_inw5;
wire [31:0] MEMOCMux48_inw6;
wire [31:0] MEMOCMux48_inw7;
wire [31:0] MEMOCMux48_inw8;
wire [31:0] MEMOCMux48_inw9;
wire [31:0] MEMOCMux48_inw10;
wire [31:0] MEMOCMux48_outw1;
wire [3:0] MEMOCMux48_selw;
HA_10IM MEMOCMux48 (
.DataIn_1(MEMOCMux48_inw1),
.DataIn_2(MEMOCMux48_inw2),
.DataIn_3(MEMOCMux48_inw3),
.DataIn_4(MEMOCMux48_inw4),
.DataIn_5(MEMOCMux48_inw5),
.DataIn_6(MEMOCMux48_inw6),
.DataIn_7(MEMOCMux48_inw7),
.DataIn_8(MEMOCMux48_inw8),
.DataIn_9(MEMOCMux48_inw9),
.DataIn_10(MEMOCMux48_inw10),
.DataOut_1(MEMOCMux48_outw1),
.sel(MEMOCMux48_selw));
defparam MEMOCMux48.Mux_BW = 32;
assign MEMC48_data_from_Core = MEMOCMux48_outw1;
assign MEMOCMux48_inw1 = dataOutW[31:0]; 
assign MEMOCMux48_inw2 = dataOutW[63:32]; 
assign MEMOCMux48_inw3 = dataOutW[95:64]; 
assign MEMOCMux48_inw4 = dataOutW[127:96]; 
assign MEMOCMux48_inw5 = dataOutW[159:128]; 
assign MEMOCMux48_inw6 = dataOutW[191:160]; 
assign MEMOCMux48_inw7 = dataOutW[223:192]; 
assign MEMOCMux48_inw8 = dataOutW[255:224]; 
assign MEMOCMux48_inw9 = dataOutW[287:256]; 
assign MEMOCMux48_inw10 = globalDataIn[1567:1536]; 
assign MEMOCMux48_selw = mOutConfigW[195:192]; 
assign MEMC48_data_out_ctx2 = mDataFromMem[1567:1536]; 
assign mDataToMem[1567:1536] = MEMC48_data_in_ctx1; 
assign globalDataOut[1567:1536] = MEMC48_data_to_Core; 
assign MEMC48_valid_ctx1 = valid1[48:48]; 
assign MEMC48_write_en_ctx1 = WEn1[48:48]; 
assign MEMC48_stride_ctx1 = stride1[48:48]; 
assign MEMC48_start_addr_ctx1 = startAddr1[293:288]; 
assign MEMC48_burst_count_ctx1 = count1[342:336]; 
assign mAddr1[293:288] = MEMC48_addr_out_ctx1; 
assign mEn1[48:48] = MEMC48_mem_en_ctx1; 
assign mWEn1[48:48] = MEMC48_write_mem_en_ctx1; 
assign MEMC48_valid_ctx2 = valid2[48:48]; 
assign MEMC48_write_en_ctx2 = WEn2[48:48]; 
assign MEMC48_stride_ctx2 = stride2[48:48]; 
assign MEMC48_start_addr_ctx2 = startAddr2[293:288]; 
assign mAddr2[293:288] = MEMC48_addr_out_ctx2; 
assign MEMC48_burst_count_ctx2 = count2[342:336]; 
assign mEn2[48:48] = MEMC48_mem_en_ctx2; 
assign mWEn2[48:48] = MEMC48_write_mem_en_ctx2; 
wire [31:0] MEMOCMux49_inw1;
wire [31:0] MEMOCMux49_inw2;
wire [31:0] MEMOCMux49_inw3;
wire [31:0] MEMOCMux49_inw4;
wire [31:0] MEMOCMux49_inw5;
wire [31:0] MEMOCMux49_inw6;
wire [31:0] MEMOCMux49_inw7;
wire [31:0] MEMOCMux49_inw8;
wire [31:0] MEMOCMux49_inw9;
wire [31:0] MEMOCMux49_inw10;
wire [31:0] MEMOCMux49_outw1;
wire [3:0] MEMOCMux49_selw;
HA_10IM MEMOCMux49 (
.DataIn_1(MEMOCMux49_inw1),
.DataIn_2(MEMOCMux49_inw2),
.DataIn_3(MEMOCMux49_inw3),
.DataIn_4(MEMOCMux49_inw4),
.DataIn_5(MEMOCMux49_inw5),
.DataIn_6(MEMOCMux49_inw6),
.DataIn_7(MEMOCMux49_inw7),
.DataIn_8(MEMOCMux49_inw8),
.DataIn_9(MEMOCMux49_inw9),
.DataIn_10(MEMOCMux49_inw10),
.DataOut_1(MEMOCMux49_outw1),
.sel(MEMOCMux49_selw));
defparam MEMOCMux49.Mux_BW = 32;
assign MEMC49_data_from_Core = MEMOCMux49_outw1;
assign MEMOCMux49_inw1 = dataOutW[31:0]; 
assign MEMOCMux49_inw2 = dataOutW[63:32]; 
assign MEMOCMux49_inw3 = dataOutW[95:64]; 
assign MEMOCMux49_inw4 = dataOutW[127:96]; 
assign MEMOCMux49_inw5 = dataOutW[159:128]; 
assign MEMOCMux49_inw6 = dataOutW[191:160]; 
assign MEMOCMux49_inw7 = dataOutW[223:192]; 
assign MEMOCMux49_inw8 = dataOutW[255:224]; 
assign MEMOCMux49_inw9 = dataOutW[287:256]; 
assign MEMOCMux49_inw10 = globalDataIn[1599:1568]; 
assign MEMOCMux49_selw = mOutConfigW[199:196]; 
assign MEMC49_data_out_ctx2 = mDataFromMem[1599:1568]; 
assign mDataToMem[1599:1568] = MEMC49_data_in_ctx1; 
assign globalDataOut[1599:1568] = MEMC49_data_to_Core; 
assign MEMC49_valid_ctx1 = valid1[49:49]; 
assign MEMC49_write_en_ctx1 = WEn1[49:49]; 
assign MEMC49_stride_ctx1 = stride1[49:49]; 
assign MEMC49_start_addr_ctx1 = startAddr1[299:294]; 
assign MEMC49_burst_count_ctx1 = count1[349:343]; 
assign mAddr1[299:294] = MEMC49_addr_out_ctx1; 
assign mEn1[49:49] = MEMC49_mem_en_ctx1; 
assign mWEn1[49:49] = MEMC49_write_mem_en_ctx1; 
assign MEMC49_valid_ctx2 = valid2[49:49]; 
assign MEMC49_write_en_ctx2 = WEn2[49:49]; 
assign MEMC49_stride_ctx2 = stride2[49:49]; 
assign MEMC49_start_addr_ctx2 = startAddr2[299:294]; 
assign mAddr2[299:294] = MEMC49_addr_out_ctx2; 
assign MEMC49_burst_count_ctx2 = count2[349:343]; 
assign mEn2[49:49] = MEMC49_mem_en_ctx2; 
assign mWEn2[49:49] = MEMC49_write_mem_en_ctx2; 
wire [31:0] MEMOCMux50_inw1;
wire [31:0] MEMOCMux50_inw2;
wire [31:0] MEMOCMux50_inw3;
wire [31:0] MEMOCMux50_inw4;
wire [31:0] MEMOCMux50_inw5;
wire [31:0] MEMOCMux50_inw6;
wire [31:0] MEMOCMux50_inw7;
wire [31:0] MEMOCMux50_inw8;
wire [31:0] MEMOCMux50_inw9;
wire [31:0] MEMOCMux50_inw10;
wire [31:0] MEMOCMux50_outw1;
wire [3:0] MEMOCMux50_selw;
HA_10IM MEMOCMux50 (
.DataIn_1(MEMOCMux50_inw1),
.DataIn_2(MEMOCMux50_inw2),
.DataIn_3(MEMOCMux50_inw3),
.DataIn_4(MEMOCMux50_inw4),
.DataIn_5(MEMOCMux50_inw5),
.DataIn_6(MEMOCMux50_inw6),
.DataIn_7(MEMOCMux50_inw7),
.DataIn_8(MEMOCMux50_inw8),
.DataIn_9(MEMOCMux50_inw9),
.DataIn_10(MEMOCMux50_inw10),
.DataOut_1(MEMOCMux50_outw1),
.sel(MEMOCMux50_selw));
defparam MEMOCMux50.Mux_BW = 32;
assign MEMC50_data_from_Core = MEMOCMux50_outw1;
assign MEMOCMux50_inw1 = dataOutW[31:0]; 
assign MEMOCMux50_inw2 = dataOutW[63:32]; 
assign MEMOCMux50_inw3 = dataOutW[95:64]; 
assign MEMOCMux50_inw4 = dataOutW[127:96]; 
assign MEMOCMux50_inw5 = dataOutW[159:128]; 
assign MEMOCMux50_inw6 = dataOutW[191:160]; 
assign MEMOCMux50_inw7 = dataOutW[223:192]; 
assign MEMOCMux50_inw8 = dataOutW[255:224]; 
assign MEMOCMux50_inw9 = dataOutW[287:256]; 
assign MEMOCMux50_inw10 = globalDataIn[1631:1600]; 
assign MEMOCMux50_selw = mOutConfigW[203:200]; 
assign MEMC50_data_out_ctx2 = mDataFromMem[1631:1600]; 
assign mDataToMem[1631:1600] = MEMC50_data_in_ctx1; 
assign globalDataOut[1631:1600] = MEMC50_data_to_Core; 
assign MEMC50_valid_ctx1 = valid1[50:50]; 
assign MEMC50_write_en_ctx1 = WEn1[50:50]; 
assign MEMC50_stride_ctx1 = stride1[50:50]; 
assign MEMC50_start_addr_ctx1 = startAddr1[305:300]; 
assign MEMC50_burst_count_ctx1 = count1[356:350]; 
assign mAddr1[305:300] = MEMC50_addr_out_ctx1; 
assign mEn1[50:50] = MEMC50_mem_en_ctx1; 
assign mWEn1[50:50] = MEMC50_write_mem_en_ctx1; 
assign MEMC50_valid_ctx2 = valid2[50:50]; 
assign MEMC50_write_en_ctx2 = WEn2[50:50]; 
assign MEMC50_stride_ctx2 = stride2[50:50]; 
assign MEMC50_start_addr_ctx2 = startAddr2[305:300]; 
assign mAddr2[305:300] = MEMC50_addr_out_ctx2; 
assign MEMC50_burst_count_ctx2 = count2[356:350]; 
assign mEn2[50:50] = MEMC50_mem_en_ctx2; 
assign mWEn2[50:50] = MEMC50_write_mem_en_ctx2; 
wire [31:0] MEMOCMux51_inw1;
wire [31:0] MEMOCMux51_inw2;
wire [31:0] MEMOCMux51_inw3;
wire [31:0] MEMOCMux51_inw4;
wire [31:0] MEMOCMux51_inw5;
wire [31:0] MEMOCMux51_inw6;
wire [31:0] MEMOCMux51_inw7;
wire [31:0] MEMOCMux51_inw8;
wire [31:0] MEMOCMux51_inw9;
wire [31:0] MEMOCMux51_inw10;
wire [31:0] MEMOCMux51_outw1;
wire [3:0] MEMOCMux51_selw;
HA_10IM MEMOCMux51 (
.DataIn_1(MEMOCMux51_inw1),
.DataIn_2(MEMOCMux51_inw2),
.DataIn_3(MEMOCMux51_inw3),
.DataIn_4(MEMOCMux51_inw4),
.DataIn_5(MEMOCMux51_inw5),
.DataIn_6(MEMOCMux51_inw6),
.DataIn_7(MEMOCMux51_inw7),
.DataIn_8(MEMOCMux51_inw8),
.DataIn_9(MEMOCMux51_inw9),
.DataIn_10(MEMOCMux51_inw10),
.DataOut_1(MEMOCMux51_outw1),
.sel(MEMOCMux51_selw));
defparam MEMOCMux51.Mux_BW = 32;
assign MEMC51_data_from_Core = MEMOCMux51_outw1;
assign MEMOCMux51_inw1 = dataOutW[31:0]; 
assign MEMOCMux51_inw2 = dataOutW[63:32]; 
assign MEMOCMux51_inw3 = dataOutW[95:64]; 
assign MEMOCMux51_inw4 = dataOutW[127:96]; 
assign MEMOCMux51_inw5 = dataOutW[159:128]; 
assign MEMOCMux51_inw6 = dataOutW[191:160]; 
assign MEMOCMux51_inw7 = dataOutW[223:192]; 
assign MEMOCMux51_inw8 = dataOutW[255:224]; 
assign MEMOCMux51_inw9 = dataOutW[287:256]; 
assign MEMOCMux51_inw10 = globalDataIn[1663:1632]; 
assign MEMOCMux51_selw = mOutConfigW[207:204]; 
assign MEMC51_data_out_ctx2 = mDataFromMem[1663:1632]; 
assign mDataToMem[1663:1632] = MEMC51_data_in_ctx1; 
assign globalDataOut[1663:1632] = MEMC51_data_to_Core; 
assign MEMC51_valid_ctx1 = valid1[51:51]; 
assign MEMC51_write_en_ctx1 = WEn1[51:51]; 
assign MEMC51_stride_ctx1 = stride1[51:51]; 
assign MEMC51_start_addr_ctx1 = startAddr1[311:306]; 
assign MEMC51_burst_count_ctx1 = count1[363:357]; 
assign mAddr1[311:306] = MEMC51_addr_out_ctx1; 
assign mEn1[51:51] = MEMC51_mem_en_ctx1; 
assign mWEn1[51:51] = MEMC51_write_mem_en_ctx1; 
assign MEMC51_valid_ctx2 = valid2[51:51]; 
assign MEMC51_write_en_ctx2 = WEn2[51:51]; 
assign MEMC51_stride_ctx2 = stride2[51:51]; 
assign MEMC51_start_addr_ctx2 = startAddr2[311:306]; 
assign mAddr2[311:306] = MEMC51_addr_out_ctx2; 
assign MEMC51_burst_count_ctx2 = count2[363:357]; 
assign mEn2[51:51] = MEMC51_mem_en_ctx2; 
assign mWEn2[51:51] = MEMC51_write_mem_en_ctx2; 
wire [31:0] MEMOCMux52_inw1;
wire [31:0] MEMOCMux52_inw2;
wire [31:0] MEMOCMux52_inw3;
wire [31:0] MEMOCMux52_inw4;
wire [31:0] MEMOCMux52_inw5;
wire [31:0] MEMOCMux52_inw6;
wire [31:0] MEMOCMux52_inw7;
wire [31:0] MEMOCMux52_inw8;
wire [31:0] MEMOCMux52_inw9;
wire [31:0] MEMOCMux52_inw10;
wire [31:0] MEMOCMux52_outw1;
wire [3:0] MEMOCMux52_selw;
HA_10IM MEMOCMux52 (
.DataIn_1(MEMOCMux52_inw1),
.DataIn_2(MEMOCMux52_inw2),
.DataIn_3(MEMOCMux52_inw3),
.DataIn_4(MEMOCMux52_inw4),
.DataIn_5(MEMOCMux52_inw5),
.DataIn_6(MEMOCMux52_inw6),
.DataIn_7(MEMOCMux52_inw7),
.DataIn_8(MEMOCMux52_inw8),
.DataIn_9(MEMOCMux52_inw9),
.DataIn_10(MEMOCMux52_inw10),
.DataOut_1(MEMOCMux52_outw1),
.sel(MEMOCMux52_selw));
defparam MEMOCMux52.Mux_BW = 32;
assign MEMC52_data_from_Core = MEMOCMux52_outw1;
assign MEMOCMux52_inw1 = dataOutW[31:0]; 
assign MEMOCMux52_inw2 = dataOutW[63:32]; 
assign MEMOCMux52_inw3 = dataOutW[95:64]; 
assign MEMOCMux52_inw4 = dataOutW[127:96]; 
assign MEMOCMux52_inw5 = dataOutW[159:128]; 
assign MEMOCMux52_inw6 = dataOutW[191:160]; 
assign MEMOCMux52_inw7 = dataOutW[223:192]; 
assign MEMOCMux52_inw8 = dataOutW[255:224]; 
assign MEMOCMux52_inw9 = dataOutW[287:256]; 
assign MEMOCMux52_inw10 = globalDataIn[1695:1664]; 
assign MEMOCMux52_selw = mOutConfigW[211:208]; 
assign MEMC52_data_out_ctx2 = mDataFromMem[1695:1664]; 
assign mDataToMem[1695:1664] = MEMC52_data_in_ctx1; 
assign globalDataOut[1695:1664] = MEMC52_data_to_Core; 
assign MEMC52_valid_ctx1 = valid1[52:52]; 
assign MEMC52_write_en_ctx1 = WEn1[52:52]; 
assign MEMC52_stride_ctx1 = stride1[52:52]; 
assign MEMC52_start_addr_ctx1 = startAddr1[317:312]; 
assign MEMC52_burst_count_ctx1 = count1[370:364]; 
assign mAddr1[317:312] = MEMC52_addr_out_ctx1; 
assign mEn1[52:52] = MEMC52_mem_en_ctx1; 
assign mWEn1[52:52] = MEMC52_write_mem_en_ctx1; 
assign MEMC52_valid_ctx2 = valid2[52:52]; 
assign MEMC52_write_en_ctx2 = WEn2[52:52]; 
assign MEMC52_stride_ctx2 = stride2[52:52]; 
assign MEMC52_start_addr_ctx2 = startAddr2[317:312]; 
assign mAddr2[317:312] = MEMC52_addr_out_ctx2; 
assign MEMC52_burst_count_ctx2 = count2[370:364]; 
assign mEn2[52:52] = MEMC52_mem_en_ctx2; 
assign mWEn2[52:52] = MEMC52_write_mem_en_ctx2; 
wire [31:0] MEMOCMux53_inw1;
wire [31:0] MEMOCMux53_inw2;
wire [31:0] MEMOCMux53_inw3;
wire [31:0] MEMOCMux53_inw4;
wire [31:0] MEMOCMux53_inw5;
wire [31:0] MEMOCMux53_inw6;
wire [31:0] MEMOCMux53_inw7;
wire [31:0] MEMOCMux53_inw8;
wire [31:0] MEMOCMux53_inw9;
wire [31:0] MEMOCMux53_inw10;
wire [31:0] MEMOCMux53_outw1;
wire [3:0] MEMOCMux53_selw;
HA_10IM MEMOCMux53 (
.DataIn_1(MEMOCMux53_inw1),
.DataIn_2(MEMOCMux53_inw2),
.DataIn_3(MEMOCMux53_inw3),
.DataIn_4(MEMOCMux53_inw4),
.DataIn_5(MEMOCMux53_inw5),
.DataIn_6(MEMOCMux53_inw6),
.DataIn_7(MEMOCMux53_inw7),
.DataIn_8(MEMOCMux53_inw8),
.DataIn_9(MEMOCMux53_inw9),
.DataIn_10(MEMOCMux53_inw10),
.DataOut_1(MEMOCMux53_outw1),
.sel(MEMOCMux53_selw));
defparam MEMOCMux53.Mux_BW = 32;
assign MEMC53_data_from_Core = MEMOCMux53_outw1;
assign MEMOCMux53_inw1 = dataOutW[31:0]; 
assign MEMOCMux53_inw2 = dataOutW[63:32]; 
assign MEMOCMux53_inw3 = dataOutW[95:64]; 
assign MEMOCMux53_inw4 = dataOutW[127:96]; 
assign MEMOCMux53_inw5 = dataOutW[159:128]; 
assign MEMOCMux53_inw6 = dataOutW[191:160]; 
assign MEMOCMux53_inw7 = dataOutW[223:192]; 
assign MEMOCMux53_inw8 = dataOutW[255:224]; 
assign MEMOCMux53_inw9 = dataOutW[287:256]; 
assign MEMOCMux53_inw10 = globalDataIn[1727:1696]; 
assign MEMOCMux53_selw = mOutConfigW[215:212]; 
assign MEMC53_data_out_ctx2 = mDataFromMem[1727:1696]; 
assign mDataToMem[1727:1696] = MEMC53_data_in_ctx1; 
assign globalDataOut[1727:1696] = MEMC53_data_to_Core; 
assign MEMC53_valid_ctx1 = valid1[53:53]; 
assign MEMC53_write_en_ctx1 = WEn1[53:53]; 
assign MEMC53_stride_ctx1 = stride1[53:53]; 
assign MEMC53_start_addr_ctx1 = startAddr1[323:318]; 
assign MEMC53_burst_count_ctx1 = count1[377:371]; 
assign mAddr1[323:318] = MEMC53_addr_out_ctx1; 
assign mEn1[53:53] = MEMC53_mem_en_ctx1; 
assign mWEn1[53:53] = MEMC53_write_mem_en_ctx1; 
assign MEMC53_valid_ctx2 = valid2[53:53]; 
assign MEMC53_write_en_ctx2 = WEn2[53:53]; 
assign MEMC53_stride_ctx2 = stride2[53:53]; 
assign MEMC53_start_addr_ctx2 = startAddr2[323:318]; 
assign mAddr2[323:318] = MEMC53_addr_out_ctx2; 
assign MEMC53_burst_count_ctx2 = count2[377:371]; 
assign mEn2[53:53] = MEMC53_mem_en_ctx2; 
assign mWEn2[53:53] = MEMC53_write_mem_en_ctx2; 
wire [31:0] MEMOCMux54_inw1;
wire [31:0] MEMOCMux54_inw2;
wire [31:0] MEMOCMux54_inw3;
wire [31:0] MEMOCMux54_inw4;
wire [31:0] MEMOCMux54_inw5;
wire [31:0] MEMOCMux54_inw6;
wire [31:0] MEMOCMux54_inw7;
wire [31:0] MEMOCMux54_inw8;
wire [31:0] MEMOCMux54_inw9;
wire [31:0] MEMOCMux54_inw10;
wire [31:0] MEMOCMux54_outw1;
wire [3:0] MEMOCMux54_selw;
HA_10IM MEMOCMux54 (
.DataIn_1(MEMOCMux54_inw1),
.DataIn_2(MEMOCMux54_inw2),
.DataIn_3(MEMOCMux54_inw3),
.DataIn_4(MEMOCMux54_inw4),
.DataIn_5(MEMOCMux54_inw5),
.DataIn_6(MEMOCMux54_inw6),
.DataIn_7(MEMOCMux54_inw7),
.DataIn_8(MEMOCMux54_inw8),
.DataIn_9(MEMOCMux54_inw9),
.DataIn_10(MEMOCMux54_inw10),
.DataOut_1(MEMOCMux54_outw1),
.sel(MEMOCMux54_selw));
defparam MEMOCMux54.Mux_BW = 32;
assign MEMC54_data_from_Core = MEMOCMux54_outw1;
assign MEMOCMux54_inw1 = dataOutW[31:0]; 
assign MEMOCMux54_inw2 = dataOutW[63:32]; 
assign MEMOCMux54_inw3 = dataOutW[95:64]; 
assign MEMOCMux54_inw4 = dataOutW[127:96]; 
assign MEMOCMux54_inw5 = dataOutW[159:128]; 
assign MEMOCMux54_inw6 = dataOutW[191:160]; 
assign MEMOCMux54_inw7 = dataOutW[223:192]; 
assign MEMOCMux54_inw8 = dataOutW[255:224]; 
assign MEMOCMux54_inw9 = dataOutW[287:256]; 
assign MEMOCMux54_inw10 = globalDataIn[1759:1728]; 
assign MEMOCMux54_selw = mOutConfigW[219:216]; 
assign MEMC54_data_out_ctx2 = mDataFromMem[1759:1728]; 
assign mDataToMem[1759:1728] = MEMC54_data_in_ctx1; 
assign globalDataOut[1759:1728] = MEMC54_data_to_Core; 
assign MEMC54_valid_ctx1 = valid1[54:54]; 
assign MEMC54_write_en_ctx1 = WEn1[54:54]; 
assign MEMC54_stride_ctx1 = stride1[54:54]; 
assign MEMC54_start_addr_ctx1 = startAddr1[329:324]; 
assign MEMC54_burst_count_ctx1 = count1[384:378]; 
assign mAddr1[329:324] = MEMC54_addr_out_ctx1; 
assign mEn1[54:54] = MEMC54_mem_en_ctx1; 
assign mWEn1[54:54] = MEMC54_write_mem_en_ctx1; 
assign MEMC54_valid_ctx2 = valid2[54:54]; 
assign MEMC54_write_en_ctx2 = WEn2[54:54]; 
assign MEMC54_stride_ctx2 = stride2[54:54]; 
assign MEMC54_start_addr_ctx2 = startAddr2[329:324]; 
assign mAddr2[329:324] = MEMC54_addr_out_ctx2; 
assign MEMC54_burst_count_ctx2 = count2[384:378]; 
assign mEn2[54:54] = MEMC54_mem_en_ctx2; 
assign mWEn2[54:54] = MEMC54_write_mem_en_ctx2; 
wire [31:0] MEMOCMux55_inw1;
wire [31:0] MEMOCMux55_inw2;
wire [31:0] MEMOCMux55_inw3;
wire [31:0] MEMOCMux55_inw4;
wire [31:0] MEMOCMux55_inw5;
wire [31:0] MEMOCMux55_inw6;
wire [31:0] MEMOCMux55_inw7;
wire [31:0] MEMOCMux55_inw8;
wire [31:0] MEMOCMux55_inw9;
wire [31:0] MEMOCMux55_inw10;
wire [31:0] MEMOCMux55_outw1;
wire [3:0] MEMOCMux55_selw;
HA_10IM MEMOCMux55 (
.DataIn_1(MEMOCMux55_inw1),
.DataIn_2(MEMOCMux55_inw2),
.DataIn_3(MEMOCMux55_inw3),
.DataIn_4(MEMOCMux55_inw4),
.DataIn_5(MEMOCMux55_inw5),
.DataIn_6(MEMOCMux55_inw6),
.DataIn_7(MEMOCMux55_inw7),
.DataIn_8(MEMOCMux55_inw8),
.DataIn_9(MEMOCMux55_inw9),
.DataIn_10(MEMOCMux55_inw10),
.DataOut_1(MEMOCMux55_outw1),
.sel(MEMOCMux55_selw));
defparam MEMOCMux55.Mux_BW = 32;
assign MEMC55_data_from_Core = MEMOCMux55_outw1;
assign MEMOCMux55_inw1 = dataOutW[31:0]; 
assign MEMOCMux55_inw2 = dataOutW[63:32]; 
assign MEMOCMux55_inw3 = dataOutW[95:64]; 
assign MEMOCMux55_inw4 = dataOutW[127:96]; 
assign MEMOCMux55_inw5 = dataOutW[159:128]; 
assign MEMOCMux55_inw6 = dataOutW[191:160]; 
assign MEMOCMux55_inw7 = dataOutW[223:192]; 
assign MEMOCMux55_inw8 = dataOutW[255:224]; 
assign MEMOCMux55_inw9 = dataOutW[287:256]; 
assign MEMOCMux55_inw10 = globalDataIn[1791:1760]; 
assign MEMOCMux55_selw = mOutConfigW[223:220]; 
assign MEMC55_data_out_ctx2 = mDataFromMem[1791:1760]; 
assign mDataToMem[1791:1760] = MEMC55_data_in_ctx1; 
assign globalDataOut[1791:1760] = MEMC55_data_to_Core; 
assign MEMC55_valid_ctx1 = valid1[55:55]; 
assign MEMC55_write_en_ctx1 = WEn1[55:55]; 
assign MEMC55_stride_ctx1 = stride1[55:55]; 
assign MEMC55_start_addr_ctx1 = startAddr1[335:330]; 
assign MEMC55_burst_count_ctx1 = count1[391:385]; 
assign mAddr1[335:330] = MEMC55_addr_out_ctx1; 
assign mEn1[55:55] = MEMC55_mem_en_ctx1; 
assign mWEn1[55:55] = MEMC55_write_mem_en_ctx1; 
assign MEMC55_valid_ctx2 = valid2[55:55]; 
assign MEMC55_write_en_ctx2 = WEn2[55:55]; 
assign MEMC55_stride_ctx2 = stride2[55:55]; 
assign MEMC55_start_addr_ctx2 = startAddr2[335:330]; 
assign mAddr2[335:330] = MEMC55_addr_out_ctx2; 
assign MEMC55_burst_count_ctx2 = count2[391:385]; 
assign mEn2[55:55] = MEMC55_mem_en_ctx2; 
assign mWEn2[55:55] = MEMC55_write_mem_en_ctx2; 
wire [31:0] MEMOCMux56_inw1;
wire [31:0] MEMOCMux56_inw2;
wire [31:0] MEMOCMux56_inw3;
wire [31:0] MEMOCMux56_inw4;
wire [31:0] MEMOCMux56_inw5;
wire [31:0] MEMOCMux56_inw6;
wire [31:0] MEMOCMux56_inw7;
wire [31:0] MEMOCMux56_inw8;
wire [31:0] MEMOCMux56_inw9;
wire [31:0] MEMOCMux56_inw10;
wire [31:0] MEMOCMux56_outw1;
wire [3:0] MEMOCMux56_selw;
HA_10IM MEMOCMux56 (
.DataIn_1(MEMOCMux56_inw1),
.DataIn_2(MEMOCMux56_inw2),
.DataIn_3(MEMOCMux56_inw3),
.DataIn_4(MEMOCMux56_inw4),
.DataIn_5(MEMOCMux56_inw5),
.DataIn_6(MEMOCMux56_inw6),
.DataIn_7(MEMOCMux56_inw7),
.DataIn_8(MEMOCMux56_inw8),
.DataIn_9(MEMOCMux56_inw9),
.DataIn_10(MEMOCMux56_inw10),
.DataOut_1(MEMOCMux56_outw1),
.sel(MEMOCMux56_selw));
defparam MEMOCMux56.Mux_BW = 32;
assign MEMC56_data_from_Core = MEMOCMux56_outw1;
assign MEMOCMux56_inw1 = dataOutW[31:0]; 
assign MEMOCMux56_inw2 = dataOutW[63:32]; 
assign MEMOCMux56_inw3 = dataOutW[95:64]; 
assign MEMOCMux56_inw4 = dataOutW[127:96]; 
assign MEMOCMux56_inw5 = dataOutW[159:128]; 
assign MEMOCMux56_inw6 = dataOutW[191:160]; 
assign MEMOCMux56_inw7 = dataOutW[223:192]; 
assign MEMOCMux56_inw8 = dataOutW[255:224]; 
assign MEMOCMux56_inw9 = dataOutW[287:256]; 
assign MEMOCMux56_inw10 = globalDataIn[1823:1792]; 
assign MEMOCMux56_selw = mOutConfigW[227:224]; 
assign MEMC56_data_out_ctx2 = mDataFromMem[1823:1792]; 
assign mDataToMem[1823:1792] = MEMC56_data_in_ctx1; 
assign globalDataOut[1823:1792] = MEMC56_data_to_Core; 
assign MEMC56_valid_ctx1 = valid1[56:56]; 
assign MEMC56_write_en_ctx1 = WEn1[56:56]; 
assign MEMC56_stride_ctx1 = stride1[56:56]; 
assign MEMC56_start_addr_ctx1 = startAddr1[341:336]; 
assign MEMC56_burst_count_ctx1 = count1[398:392]; 
assign mAddr1[341:336] = MEMC56_addr_out_ctx1; 
assign mEn1[56:56] = MEMC56_mem_en_ctx1; 
assign mWEn1[56:56] = MEMC56_write_mem_en_ctx1; 
assign MEMC56_valid_ctx2 = valid2[56:56]; 
assign MEMC56_write_en_ctx2 = WEn2[56:56]; 
assign MEMC56_stride_ctx2 = stride2[56:56]; 
assign MEMC56_start_addr_ctx2 = startAddr2[341:336]; 
assign mAddr2[341:336] = MEMC56_addr_out_ctx2; 
assign MEMC56_burst_count_ctx2 = count2[398:392]; 
assign mEn2[56:56] = MEMC56_mem_en_ctx2; 
assign mWEn2[56:56] = MEMC56_write_mem_en_ctx2; 
wire [31:0] MEMOCMux57_inw1;
wire [31:0] MEMOCMux57_inw2;
wire [31:0] MEMOCMux57_inw3;
wire [31:0] MEMOCMux57_inw4;
wire [31:0] MEMOCMux57_inw5;
wire [31:0] MEMOCMux57_inw6;
wire [31:0] MEMOCMux57_inw7;
wire [31:0] MEMOCMux57_inw8;
wire [31:0] MEMOCMux57_inw9;
wire [31:0] MEMOCMux57_inw10;
wire [31:0] MEMOCMux57_outw1;
wire [3:0] MEMOCMux57_selw;
HA_10IM MEMOCMux57 (
.DataIn_1(MEMOCMux57_inw1),
.DataIn_2(MEMOCMux57_inw2),
.DataIn_3(MEMOCMux57_inw3),
.DataIn_4(MEMOCMux57_inw4),
.DataIn_5(MEMOCMux57_inw5),
.DataIn_6(MEMOCMux57_inw6),
.DataIn_7(MEMOCMux57_inw7),
.DataIn_8(MEMOCMux57_inw8),
.DataIn_9(MEMOCMux57_inw9),
.DataIn_10(MEMOCMux57_inw10),
.DataOut_1(MEMOCMux57_outw1),
.sel(MEMOCMux57_selw));
defparam MEMOCMux57.Mux_BW = 32;
assign MEMC57_data_from_Core = MEMOCMux57_outw1;
assign MEMOCMux57_inw1 = dataOutW[31:0]; 
assign MEMOCMux57_inw2 = dataOutW[63:32]; 
assign MEMOCMux57_inw3 = dataOutW[95:64]; 
assign MEMOCMux57_inw4 = dataOutW[127:96]; 
assign MEMOCMux57_inw5 = dataOutW[159:128]; 
assign MEMOCMux57_inw6 = dataOutW[191:160]; 
assign MEMOCMux57_inw7 = dataOutW[223:192]; 
assign MEMOCMux57_inw8 = dataOutW[255:224]; 
assign MEMOCMux57_inw9 = dataOutW[287:256]; 
assign MEMOCMux57_inw10 = globalDataIn[1855:1824]; 
assign MEMOCMux57_selw = mOutConfigW[231:228]; 
assign MEMC57_data_out_ctx2 = mDataFromMem[1855:1824]; 
assign mDataToMem[1855:1824] = MEMC57_data_in_ctx1; 
assign globalDataOut[1855:1824] = MEMC57_data_to_Core; 
assign MEMC57_valid_ctx1 = valid1[57:57]; 
assign MEMC57_write_en_ctx1 = WEn1[57:57]; 
assign MEMC57_stride_ctx1 = stride1[57:57]; 
assign MEMC57_start_addr_ctx1 = startAddr1[347:342]; 
assign MEMC57_burst_count_ctx1 = count1[405:399]; 
assign mAddr1[347:342] = MEMC57_addr_out_ctx1; 
assign mEn1[57:57] = MEMC57_mem_en_ctx1; 
assign mWEn1[57:57] = MEMC57_write_mem_en_ctx1; 
assign MEMC57_valid_ctx2 = valid2[57:57]; 
assign MEMC57_write_en_ctx2 = WEn2[57:57]; 
assign MEMC57_stride_ctx2 = stride2[57:57]; 
assign MEMC57_start_addr_ctx2 = startAddr2[347:342]; 
assign mAddr2[347:342] = MEMC57_addr_out_ctx2; 
assign MEMC57_burst_count_ctx2 = count2[405:399]; 
assign mEn2[57:57] = MEMC57_mem_en_ctx2; 
assign mWEn2[57:57] = MEMC57_write_mem_en_ctx2; 
wire [31:0] MEMOCMux58_inw1;
wire [31:0] MEMOCMux58_inw2;
wire [31:0] MEMOCMux58_inw3;
wire [31:0] MEMOCMux58_inw4;
wire [31:0] MEMOCMux58_inw5;
wire [31:0] MEMOCMux58_inw6;
wire [31:0] MEMOCMux58_inw7;
wire [31:0] MEMOCMux58_inw8;
wire [31:0] MEMOCMux58_inw9;
wire [31:0] MEMOCMux58_inw10;
wire [31:0] MEMOCMux58_outw1;
wire [3:0] MEMOCMux58_selw;
HA_10IM MEMOCMux58 (
.DataIn_1(MEMOCMux58_inw1),
.DataIn_2(MEMOCMux58_inw2),
.DataIn_3(MEMOCMux58_inw3),
.DataIn_4(MEMOCMux58_inw4),
.DataIn_5(MEMOCMux58_inw5),
.DataIn_6(MEMOCMux58_inw6),
.DataIn_7(MEMOCMux58_inw7),
.DataIn_8(MEMOCMux58_inw8),
.DataIn_9(MEMOCMux58_inw9),
.DataIn_10(MEMOCMux58_inw10),
.DataOut_1(MEMOCMux58_outw1),
.sel(MEMOCMux58_selw));
defparam MEMOCMux58.Mux_BW = 32;
assign MEMC58_data_from_Core = MEMOCMux58_outw1;
assign MEMOCMux58_inw1 = dataOutW[31:0]; 
assign MEMOCMux58_inw2 = dataOutW[63:32]; 
assign MEMOCMux58_inw3 = dataOutW[95:64]; 
assign MEMOCMux58_inw4 = dataOutW[127:96]; 
assign MEMOCMux58_inw5 = dataOutW[159:128]; 
assign MEMOCMux58_inw6 = dataOutW[191:160]; 
assign MEMOCMux58_inw7 = dataOutW[223:192]; 
assign MEMOCMux58_inw8 = dataOutW[255:224]; 
assign MEMOCMux58_inw9 = dataOutW[287:256]; 
assign MEMOCMux58_inw10 = globalDataIn[1887:1856]; 
assign MEMOCMux58_selw = mOutConfigW[235:232]; 
assign MEMC58_data_out_ctx2 = mDataFromMem[1887:1856]; 
assign mDataToMem[1887:1856] = MEMC58_data_in_ctx1; 
assign globalDataOut[1887:1856] = MEMC58_data_to_Core; 
assign MEMC58_valid_ctx1 = valid1[58:58]; 
assign MEMC58_write_en_ctx1 = WEn1[58:58]; 
assign MEMC58_stride_ctx1 = stride1[58:58]; 
assign MEMC58_start_addr_ctx1 = startAddr1[353:348]; 
assign MEMC58_burst_count_ctx1 = count1[412:406]; 
assign mAddr1[353:348] = MEMC58_addr_out_ctx1; 
assign mEn1[58:58] = MEMC58_mem_en_ctx1; 
assign mWEn1[58:58] = MEMC58_write_mem_en_ctx1; 
assign MEMC58_valid_ctx2 = valid2[58:58]; 
assign MEMC58_write_en_ctx2 = WEn2[58:58]; 
assign MEMC58_stride_ctx2 = stride2[58:58]; 
assign MEMC58_start_addr_ctx2 = startAddr2[353:348]; 
assign mAddr2[353:348] = MEMC58_addr_out_ctx2; 
assign MEMC58_burst_count_ctx2 = count2[412:406]; 
assign mEn2[58:58] = MEMC58_mem_en_ctx2; 
assign mWEn2[58:58] = MEMC58_write_mem_en_ctx2; 
wire [31:0] MEMOCMux59_inw1;
wire [31:0] MEMOCMux59_inw2;
wire [31:0] MEMOCMux59_inw3;
wire [31:0] MEMOCMux59_inw4;
wire [31:0] MEMOCMux59_inw5;
wire [31:0] MEMOCMux59_inw6;
wire [31:0] MEMOCMux59_inw7;
wire [31:0] MEMOCMux59_inw8;
wire [31:0] MEMOCMux59_inw9;
wire [31:0] MEMOCMux59_inw10;
wire [31:0] MEMOCMux59_outw1;
wire [3:0] MEMOCMux59_selw;
HA_10IM MEMOCMux59 (
.DataIn_1(MEMOCMux59_inw1),
.DataIn_2(MEMOCMux59_inw2),
.DataIn_3(MEMOCMux59_inw3),
.DataIn_4(MEMOCMux59_inw4),
.DataIn_5(MEMOCMux59_inw5),
.DataIn_6(MEMOCMux59_inw6),
.DataIn_7(MEMOCMux59_inw7),
.DataIn_8(MEMOCMux59_inw8),
.DataIn_9(MEMOCMux59_inw9),
.DataIn_10(MEMOCMux59_inw10),
.DataOut_1(MEMOCMux59_outw1),
.sel(MEMOCMux59_selw));
defparam MEMOCMux59.Mux_BW = 32;
assign MEMC59_data_from_Core = MEMOCMux59_outw1;
assign MEMOCMux59_inw1 = dataOutW[31:0]; 
assign MEMOCMux59_inw2 = dataOutW[63:32]; 
assign MEMOCMux59_inw3 = dataOutW[95:64]; 
assign MEMOCMux59_inw4 = dataOutW[127:96]; 
assign MEMOCMux59_inw5 = dataOutW[159:128]; 
assign MEMOCMux59_inw6 = dataOutW[191:160]; 
assign MEMOCMux59_inw7 = dataOutW[223:192]; 
assign MEMOCMux59_inw8 = dataOutW[255:224]; 
assign MEMOCMux59_inw9 = dataOutW[287:256]; 
assign MEMOCMux59_inw10 = globalDataIn[1919:1888]; 
assign MEMOCMux59_selw = mOutConfigW[239:236]; 
assign MEMC59_data_out_ctx2 = mDataFromMem[1919:1888]; 
assign mDataToMem[1919:1888] = MEMC59_data_in_ctx1; 
assign globalDataOut[1919:1888] = MEMC59_data_to_Core; 
assign MEMC59_valid_ctx1 = valid1[59:59]; 
assign MEMC59_write_en_ctx1 = WEn1[59:59]; 
assign MEMC59_stride_ctx1 = stride1[59:59]; 
assign MEMC59_start_addr_ctx1 = startAddr1[359:354]; 
assign MEMC59_burst_count_ctx1 = count1[419:413]; 
assign mAddr1[359:354] = MEMC59_addr_out_ctx1; 
assign mEn1[59:59] = MEMC59_mem_en_ctx1; 
assign mWEn1[59:59] = MEMC59_write_mem_en_ctx1; 
assign MEMC59_valid_ctx2 = valid2[59:59]; 
assign MEMC59_write_en_ctx2 = WEn2[59:59]; 
assign MEMC59_stride_ctx2 = stride2[59:59]; 
assign MEMC59_start_addr_ctx2 = startAddr2[359:354]; 
assign mAddr2[359:354] = MEMC59_addr_out_ctx2; 
assign MEMC59_burst_count_ctx2 = count2[419:413]; 
assign mEn2[59:59] = MEMC59_mem_en_ctx2; 
assign mWEn2[59:59] = MEMC59_write_mem_en_ctx2; 
wire [31:0] MEMOCMux60_inw1;
wire [31:0] MEMOCMux60_inw2;
wire [31:0] MEMOCMux60_inw3;
wire [31:0] MEMOCMux60_inw4;
wire [31:0] MEMOCMux60_inw5;
wire [31:0] MEMOCMux60_inw6;
wire [31:0] MEMOCMux60_inw7;
wire [31:0] MEMOCMux60_inw8;
wire [31:0] MEMOCMux60_inw9;
wire [31:0] MEMOCMux60_inw10;
wire [31:0] MEMOCMux60_outw1;
wire [3:0] MEMOCMux60_selw;
HA_10IM MEMOCMux60 (
.DataIn_1(MEMOCMux60_inw1),
.DataIn_2(MEMOCMux60_inw2),
.DataIn_3(MEMOCMux60_inw3),
.DataIn_4(MEMOCMux60_inw4),
.DataIn_5(MEMOCMux60_inw5),
.DataIn_6(MEMOCMux60_inw6),
.DataIn_7(MEMOCMux60_inw7),
.DataIn_8(MEMOCMux60_inw8),
.DataIn_9(MEMOCMux60_inw9),
.DataIn_10(MEMOCMux60_inw10),
.DataOut_1(MEMOCMux60_outw1),
.sel(MEMOCMux60_selw));
defparam MEMOCMux60.Mux_BW = 32;
assign MEMC60_data_from_Core = MEMOCMux60_outw1;
assign MEMOCMux60_inw1 = dataOutW[31:0]; 
assign MEMOCMux60_inw2 = dataOutW[63:32]; 
assign MEMOCMux60_inw3 = dataOutW[95:64]; 
assign MEMOCMux60_inw4 = dataOutW[127:96]; 
assign MEMOCMux60_inw5 = dataOutW[159:128]; 
assign MEMOCMux60_inw6 = dataOutW[191:160]; 
assign MEMOCMux60_inw7 = dataOutW[223:192]; 
assign MEMOCMux60_inw8 = dataOutW[255:224]; 
assign MEMOCMux60_inw9 = dataOutW[287:256]; 
assign MEMOCMux60_inw10 = globalDataIn[1951:1920]; 
assign MEMOCMux60_selw = mOutConfigW[243:240]; 
assign MEMC60_data_out_ctx2 = mDataFromMem[1951:1920]; 
assign mDataToMem[1951:1920] = MEMC60_data_in_ctx1; 
assign globalDataOut[1951:1920] = MEMC60_data_to_Core; 
assign MEMC60_valid_ctx1 = valid1[60:60]; 
assign MEMC60_write_en_ctx1 = WEn1[60:60]; 
assign MEMC60_stride_ctx1 = stride1[60:60]; 
assign MEMC60_start_addr_ctx1 = startAddr1[365:360]; 
assign MEMC60_burst_count_ctx1 = count1[426:420]; 
assign mAddr1[365:360] = MEMC60_addr_out_ctx1; 
assign mEn1[60:60] = MEMC60_mem_en_ctx1; 
assign mWEn1[60:60] = MEMC60_write_mem_en_ctx1; 
assign MEMC60_valid_ctx2 = valid2[60:60]; 
assign MEMC60_write_en_ctx2 = WEn2[60:60]; 
assign MEMC60_stride_ctx2 = stride2[60:60]; 
assign MEMC60_start_addr_ctx2 = startAddr2[365:360]; 
assign mAddr2[365:360] = MEMC60_addr_out_ctx2; 
assign MEMC60_burst_count_ctx2 = count2[426:420]; 
assign mEn2[60:60] = MEMC60_mem_en_ctx2; 
assign mWEn2[60:60] = MEMC60_write_mem_en_ctx2; 
wire [31:0] MEMOCMux61_inw1;
wire [31:0] MEMOCMux61_inw2;
wire [31:0] MEMOCMux61_inw3;
wire [31:0] MEMOCMux61_inw4;
wire [31:0] MEMOCMux61_inw5;
wire [31:0] MEMOCMux61_inw6;
wire [31:0] MEMOCMux61_inw7;
wire [31:0] MEMOCMux61_inw8;
wire [31:0] MEMOCMux61_inw9;
wire [31:0] MEMOCMux61_inw10;
wire [31:0] MEMOCMux61_outw1;
wire [3:0] MEMOCMux61_selw;
HA_10IM MEMOCMux61 (
.DataIn_1(MEMOCMux61_inw1),
.DataIn_2(MEMOCMux61_inw2),
.DataIn_3(MEMOCMux61_inw3),
.DataIn_4(MEMOCMux61_inw4),
.DataIn_5(MEMOCMux61_inw5),
.DataIn_6(MEMOCMux61_inw6),
.DataIn_7(MEMOCMux61_inw7),
.DataIn_8(MEMOCMux61_inw8),
.DataIn_9(MEMOCMux61_inw9),
.DataIn_10(MEMOCMux61_inw10),
.DataOut_1(MEMOCMux61_outw1),
.sel(MEMOCMux61_selw));
defparam MEMOCMux61.Mux_BW = 32;
assign MEMC61_data_from_Core = MEMOCMux61_outw1;
assign MEMOCMux61_inw1 = dataOutW[31:0]; 
assign MEMOCMux61_inw2 = dataOutW[63:32]; 
assign MEMOCMux61_inw3 = dataOutW[95:64]; 
assign MEMOCMux61_inw4 = dataOutW[127:96]; 
assign MEMOCMux61_inw5 = dataOutW[159:128]; 
assign MEMOCMux61_inw6 = dataOutW[191:160]; 
assign MEMOCMux61_inw7 = dataOutW[223:192]; 
assign MEMOCMux61_inw8 = dataOutW[255:224]; 
assign MEMOCMux61_inw9 = dataOutW[287:256]; 
assign MEMOCMux61_inw10 = globalDataIn[1983:1952]; 
assign MEMOCMux61_selw = mOutConfigW[247:244]; 
assign MEMC61_data_out_ctx2 = mDataFromMem[1983:1952]; 
assign mDataToMem[1983:1952] = MEMC61_data_in_ctx1; 
assign globalDataOut[1983:1952] = MEMC61_data_to_Core; 
assign MEMC61_valid_ctx1 = valid1[61:61]; 
assign MEMC61_write_en_ctx1 = WEn1[61:61]; 
assign MEMC61_stride_ctx1 = stride1[61:61]; 
assign MEMC61_start_addr_ctx1 = startAddr1[371:366]; 
assign MEMC61_burst_count_ctx1 = count1[433:427]; 
assign mAddr1[371:366] = MEMC61_addr_out_ctx1; 
assign mEn1[61:61] = MEMC61_mem_en_ctx1; 
assign mWEn1[61:61] = MEMC61_write_mem_en_ctx1; 
assign MEMC61_valid_ctx2 = valid2[61:61]; 
assign MEMC61_write_en_ctx2 = WEn2[61:61]; 
assign MEMC61_stride_ctx2 = stride2[61:61]; 
assign MEMC61_start_addr_ctx2 = startAddr2[371:366]; 
assign mAddr2[371:366] = MEMC61_addr_out_ctx2; 
assign MEMC61_burst_count_ctx2 = count2[433:427]; 
assign mEn2[61:61] = MEMC61_mem_en_ctx2; 
assign mWEn2[61:61] = MEMC61_write_mem_en_ctx2; 
wire [31:0] MEMOCMux62_inw1;
wire [31:0] MEMOCMux62_inw2;
wire [31:0] MEMOCMux62_inw3;
wire [31:0] MEMOCMux62_inw4;
wire [31:0] MEMOCMux62_inw5;
wire [31:0] MEMOCMux62_inw6;
wire [31:0] MEMOCMux62_inw7;
wire [31:0] MEMOCMux62_inw8;
wire [31:0] MEMOCMux62_inw9;
wire [31:0] MEMOCMux62_inw10;
wire [31:0] MEMOCMux62_outw1;
wire [3:0] MEMOCMux62_selw;
HA_10IM MEMOCMux62 (
.DataIn_1(MEMOCMux62_inw1),
.DataIn_2(MEMOCMux62_inw2),
.DataIn_3(MEMOCMux62_inw3),
.DataIn_4(MEMOCMux62_inw4),
.DataIn_5(MEMOCMux62_inw5),
.DataIn_6(MEMOCMux62_inw6),
.DataIn_7(MEMOCMux62_inw7),
.DataIn_8(MEMOCMux62_inw8),
.DataIn_9(MEMOCMux62_inw9),
.DataIn_10(MEMOCMux62_inw10),
.DataOut_1(MEMOCMux62_outw1),
.sel(MEMOCMux62_selw));
defparam MEMOCMux62.Mux_BW = 32;
assign MEMC62_data_from_Core = MEMOCMux62_outw1;
assign MEMOCMux62_inw1 = dataOutW[31:0]; 
assign MEMOCMux62_inw2 = dataOutW[63:32]; 
assign MEMOCMux62_inw3 = dataOutW[95:64]; 
assign MEMOCMux62_inw4 = dataOutW[127:96]; 
assign MEMOCMux62_inw5 = dataOutW[159:128]; 
assign MEMOCMux62_inw6 = dataOutW[191:160]; 
assign MEMOCMux62_inw7 = dataOutW[223:192]; 
assign MEMOCMux62_inw8 = dataOutW[255:224]; 
assign MEMOCMux62_inw9 = dataOutW[287:256]; 
assign MEMOCMux62_inw10 = globalDataIn[2015:1984]; 
assign MEMOCMux62_selw = mOutConfigW[251:248]; 
assign MEMC62_data_out_ctx2 = mDataFromMem[2015:1984]; 
assign mDataToMem[2015:1984] = MEMC62_data_in_ctx1; 
assign globalDataOut[2015:1984] = MEMC62_data_to_Core; 
assign MEMC62_valid_ctx1 = valid1[62:62]; 
assign MEMC62_write_en_ctx1 = WEn1[62:62]; 
assign MEMC62_stride_ctx1 = stride1[62:62]; 
assign MEMC62_start_addr_ctx1 = startAddr1[377:372]; 
assign MEMC62_burst_count_ctx1 = count1[440:434]; 
assign mAddr1[377:372] = MEMC62_addr_out_ctx1; 
assign mEn1[62:62] = MEMC62_mem_en_ctx1; 
assign mWEn1[62:62] = MEMC62_write_mem_en_ctx1; 
assign MEMC62_valid_ctx2 = valid2[62:62]; 
assign MEMC62_write_en_ctx2 = WEn2[62:62]; 
assign MEMC62_stride_ctx2 = stride2[62:62]; 
assign MEMC62_start_addr_ctx2 = startAddr2[377:372]; 
assign mAddr2[377:372] = MEMC62_addr_out_ctx2; 
assign MEMC62_burst_count_ctx2 = count2[440:434]; 
assign mEn2[62:62] = MEMC62_mem_en_ctx2; 
assign mWEn2[62:62] = MEMC62_write_mem_en_ctx2; 
wire [31:0] MEMOCMux63_inw1;
wire [31:0] MEMOCMux63_inw2;
wire [31:0] MEMOCMux63_inw3;
wire [31:0] MEMOCMux63_inw4;
wire [31:0] MEMOCMux63_inw5;
wire [31:0] MEMOCMux63_inw6;
wire [31:0] MEMOCMux63_inw7;
wire [31:0] MEMOCMux63_inw8;
wire [31:0] MEMOCMux63_inw9;
wire [31:0] MEMOCMux63_inw10;
wire [31:0] MEMOCMux63_outw1;
wire [3:0] MEMOCMux63_selw;
HA_10IM MEMOCMux63 (
.DataIn_1(MEMOCMux63_inw1),
.DataIn_2(MEMOCMux63_inw2),
.DataIn_3(MEMOCMux63_inw3),
.DataIn_4(MEMOCMux63_inw4),
.DataIn_5(MEMOCMux63_inw5),
.DataIn_6(MEMOCMux63_inw6),
.DataIn_7(MEMOCMux63_inw7),
.DataIn_8(MEMOCMux63_inw8),
.DataIn_9(MEMOCMux63_inw9),
.DataIn_10(MEMOCMux63_inw10),
.DataOut_1(MEMOCMux63_outw1),
.sel(MEMOCMux63_selw));
defparam MEMOCMux63.Mux_BW = 32;
assign MEMC63_data_from_Core = MEMOCMux63_outw1;
assign MEMOCMux63_inw1 = dataOutW[31:0]; 
assign MEMOCMux63_inw2 = dataOutW[63:32]; 
assign MEMOCMux63_inw3 = dataOutW[95:64]; 
assign MEMOCMux63_inw4 = dataOutW[127:96]; 
assign MEMOCMux63_inw5 = dataOutW[159:128]; 
assign MEMOCMux63_inw6 = dataOutW[191:160]; 
assign MEMOCMux63_inw7 = dataOutW[223:192]; 
assign MEMOCMux63_inw8 = dataOutW[255:224]; 
assign MEMOCMux63_inw9 = dataOutW[287:256]; 
assign MEMOCMux63_inw10 = globalDataIn[2047:2016]; 
assign MEMOCMux63_selw = mOutConfigW[255:252]; 
assign MEMC63_data_out_ctx2 = mDataFromMem[2047:2016]; 
assign mDataToMem[2047:2016] = MEMC63_data_in_ctx1; 
assign globalDataOut[2047:2016] = MEMC63_data_to_Core; 
assign MEMC63_valid_ctx1 = valid1[63:63]; 
assign MEMC63_write_en_ctx1 = WEn1[63:63]; 
assign MEMC63_stride_ctx1 = stride1[63:63]; 
assign MEMC63_start_addr_ctx1 = startAddr1[383:378]; 
assign MEMC63_burst_count_ctx1 = count1[447:441]; 
assign mAddr1[383:378] = MEMC63_addr_out_ctx1; 
assign mEn1[63:63] = MEMC63_mem_en_ctx1; 
assign mWEn1[63:63] = MEMC63_write_mem_en_ctx1; 
assign MEMC63_valid_ctx2 = valid2[63:63]; 
assign MEMC63_write_en_ctx2 = WEn2[63:63]; 
assign MEMC63_stride_ctx2 = stride2[63:63]; 
assign MEMC63_start_addr_ctx2 = startAddr2[383:378]; 
assign mAddr2[383:378] = MEMC63_addr_out_ctx2; 
assign MEMC63_burst_count_ctx2 = count2[447:441]; 
assign mEn2[63:63] = MEMC63_mem_en_ctx2; 
assign mWEn2[63:63] = MEMC63_write_mem_en_ctx2; 
wire [31:0] MEMOCMux64_inw1;
wire [31:0] MEMOCMux64_inw2;
wire [31:0] MEMOCMux64_inw3;
wire [31:0] MEMOCMux64_inw4;
wire [31:0] MEMOCMux64_inw5;
wire [31:0] MEMOCMux64_inw6;
wire [31:0] MEMOCMux64_inw7;
wire [31:0] MEMOCMux64_inw8;
wire [31:0] MEMOCMux64_inw9;
wire [31:0] MEMOCMux64_inw10;
wire [31:0] MEMOCMux64_outw1;
wire [3:0] MEMOCMux64_selw;
HA_10IM MEMOCMux64 (
.DataIn_1(MEMOCMux64_inw1),
.DataIn_2(MEMOCMux64_inw2),
.DataIn_3(MEMOCMux64_inw3),
.DataIn_4(MEMOCMux64_inw4),
.DataIn_5(MEMOCMux64_inw5),
.DataIn_6(MEMOCMux64_inw6),
.DataIn_7(MEMOCMux64_inw7),
.DataIn_8(MEMOCMux64_inw8),
.DataIn_9(MEMOCMux64_inw9),
.DataIn_10(MEMOCMux64_inw10),
.DataOut_1(MEMOCMux64_outw1),
.sel(MEMOCMux64_selw));
defparam MEMOCMux64.Mux_BW = 32;
assign MEMC64_data_from_Core = MEMOCMux64_outw1;
assign MEMOCMux64_inw1 = dataOutW[31:0]; 
assign MEMOCMux64_inw2 = dataOutW[63:32]; 
assign MEMOCMux64_inw3 = dataOutW[95:64]; 
assign MEMOCMux64_inw4 = dataOutW[127:96]; 
assign MEMOCMux64_inw5 = dataOutW[159:128]; 
assign MEMOCMux64_inw6 = dataOutW[191:160]; 
assign MEMOCMux64_inw7 = dataOutW[223:192]; 
assign MEMOCMux64_inw8 = dataOutW[255:224]; 
assign MEMOCMux64_inw9 = dataOutW[287:256]; 
assign MEMOCMux64_inw10 = globalDataIn[2079:2048]; 
assign MEMOCMux64_selw = mOutConfigW[259:256]; 
assign MEMC64_data_out_ctx2 = mDataFromMem[2079:2048]; 
assign mDataToMem[2079:2048] = MEMC64_data_in_ctx1; 
assign globalDataOut[2079:2048] = MEMC64_data_to_Core; 
assign MEMC64_valid_ctx1 = valid1[64:64]; 
assign MEMC64_write_en_ctx1 = WEn1[64:64]; 
assign MEMC64_stride_ctx1 = stride1[64:64]; 
assign MEMC64_start_addr_ctx1 = startAddr1[389:384]; 
assign MEMC64_burst_count_ctx1 = count1[454:448]; 
assign mAddr1[389:384] = MEMC64_addr_out_ctx1; 
assign mEn1[64:64] = MEMC64_mem_en_ctx1; 
assign mWEn1[64:64] = MEMC64_write_mem_en_ctx1; 
assign MEMC64_valid_ctx2 = valid2[64:64]; 
assign MEMC64_write_en_ctx2 = WEn2[64:64]; 
assign MEMC64_stride_ctx2 = stride2[64:64]; 
assign MEMC64_start_addr_ctx2 = startAddr2[389:384]; 
assign mAddr2[389:384] = MEMC64_addr_out_ctx2; 
assign MEMC64_burst_count_ctx2 = count2[454:448]; 
assign mEn2[64:64] = MEMC64_mem_en_ctx2; 
assign mWEn2[64:64] = MEMC64_write_mem_en_ctx2; 
wire [31:0] MEMOCMux65_inw1;
wire [31:0] MEMOCMux65_inw2;
wire [31:0] MEMOCMux65_inw3;
wire [31:0] MEMOCMux65_inw4;
wire [31:0] MEMOCMux65_inw5;
wire [31:0] MEMOCMux65_inw6;
wire [31:0] MEMOCMux65_inw7;
wire [31:0] MEMOCMux65_inw8;
wire [31:0] MEMOCMux65_inw9;
wire [31:0] MEMOCMux65_inw10;
wire [31:0] MEMOCMux65_outw1;
wire [3:0] MEMOCMux65_selw;
HA_10IM MEMOCMux65 (
.DataIn_1(MEMOCMux65_inw1),
.DataIn_2(MEMOCMux65_inw2),
.DataIn_3(MEMOCMux65_inw3),
.DataIn_4(MEMOCMux65_inw4),
.DataIn_5(MEMOCMux65_inw5),
.DataIn_6(MEMOCMux65_inw6),
.DataIn_7(MEMOCMux65_inw7),
.DataIn_8(MEMOCMux65_inw8),
.DataIn_9(MEMOCMux65_inw9),
.DataIn_10(MEMOCMux65_inw10),
.DataOut_1(MEMOCMux65_outw1),
.sel(MEMOCMux65_selw));
defparam MEMOCMux65.Mux_BW = 32;
assign MEMC65_data_from_Core = MEMOCMux65_outw1;
assign MEMOCMux65_inw1 = dataOutW[31:0]; 
assign MEMOCMux65_inw2 = dataOutW[63:32]; 
assign MEMOCMux65_inw3 = dataOutW[95:64]; 
assign MEMOCMux65_inw4 = dataOutW[127:96]; 
assign MEMOCMux65_inw5 = dataOutW[159:128]; 
assign MEMOCMux65_inw6 = dataOutW[191:160]; 
assign MEMOCMux65_inw7 = dataOutW[223:192]; 
assign MEMOCMux65_inw8 = dataOutW[255:224]; 
assign MEMOCMux65_inw9 = dataOutW[287:256]; 
assign MEMOCMux65_inw10 = globalDataIn[2111:2080]; 
assign MEMOCMux65_selw = mOutConfigW[263:260]; 
assign MEMC65_data_out_ctx2 = mDataFromMem[2111:2080]; 
assign mDataToMem[2111:2080] = MEMC65_data_in_ctx1; 
assign globalDataOut[2111:2080] = MEMC65_data_to_Core; 
assign MEMC65_valid_ctx1 = valid1[65:65]; 
assign MEMC65_write_en_ctx1 = WEn1[65:65]; 
assign MEMC65_stride_ctx1 = stride1[65:65]; 
assign MEMC65_start_addr_ctx1 = startAddr1[395:390]; 
assign MEMC65_burst_count_ctx1 = count1[461:455]; 
assign mAddr1[395:390] = MEMC65_addr_out_ctx1; 
assign mEn1[65:65] = MEMC65_mem_en_ctx1; 
assign mWEn1[65:65] = MEMC65_write_mem_en_ctx1; 
assign MEMC65_valid_ctx2 = valid2[65:65]; 
assign MEMC65_write_en_ctx2 = WEn2[65:65]; 
assign MEMC65_stride_ctx2 = stride2[65:65]; 
assign MEMC65_start_addr_ctx2 = startAddr2[395:390]; 
assign mAddr2[395:390] = MEMC65_addr_out_ctx2; 
assign MEMC65_burst_count_ctx2 = count2[461:455]; 
assign mEn2[65:65] = MEMC65_mem_en_ctx2; 
assign mWEn2[65:65] = MEMC65_write_mem_en_ctx2; 
wire [31:0] MEMOCMux66_inw1;
wire [31:0] MEMOCMux66_inw2;
wire [31:0] MEMOCMux66_inw3;
wire [31:0] MEMOCMux66_inw4;
wire [31:0] MEMOCMux66_inw5;
wire [31:0] MEMOCMux66_inw6;
wire [31:0] MEMOCMux66_inw7;
wire [31:0] MEMOCMux66_inw8;
wire [31:0] MEMOCMux66_inw9;
wire [31:0] MEMOCMux66_inw10;
wire [31:0] MEMOCMux66_outw1;
wire [3:0] MEMOCMux66_selw;
HA_10IM MEMOCMux66 (
.DataIn_1(MEMOCMux66_inw1),
.DataIn_2(MEMOCMux66_inw2),
.DataIn_3(MEMOCMux66_inw3),
.DataIn_4(MEMOCMux66_inw4),
.DataIn_5(MEMOCMux66_inw5),
.DataIn_6(MEMOCMux66_inw6),
.DataIn_7(MEMOCMux66_inw7),
.DataIn_8(MEMOCMux66_inw8),
.DataIn_9(MEMOCMux66_inw9),
.DataIn_10(MEMOCMux66_inw10),
.DataOut_1(MEMOCMux66_outw1),
.sel(MEMOCMux66_selw));
defparam MEMOCMux66.Mux_BW = 32;
assign MEMC66_data_from_Core = MEMOCMux66_outw1;
assign MEMOCMux66_inw1 = dataOutW[31:0]; 
assign MEMOCMux66_inw2 = dataOutW[63:32]; 
assign MEMOCMux66_inw3 = dataOutW[95:64]; 
assign MEMOCMux66_inw4 = dataOutW[127:96]; 
assign MEMOCMux66_inw5 = dataOutW[159:128]; 
assign MEMOCMux66_inw6 = dataOutW[191:160]; 
assign MEMOCMux66_inw7 = dataOutW[223:192]; 
assign MEMOCMux66_inw8 = dataOutW[255:224]; 
assign MEMOCMux66_inw9 = dataOutW[287:256]; 
assign MEMOCMux66_inw10 = globalDataIn[2143:2112]; 
assign MEMOCMux66_selw = mOutConfigW[267:264]; 
assign MEMC66_data_out_ctx2 = mDataFromMem[2143:2112]; 
assign mDataToMem[2143:2112] = MEMC66_data_in_ctx1; 
assign globalDataOut[2143:2112] = MEMC66_data_to_Core; 
assign MEMC66_valid_ctx1 = valid1[66:66]; 
assign MEMC66_write_en_ctx1 = WEn1[66:66]; 
assign MEMC66_stride_ctx1 = stride1[66:66]; 
assign MEMC66_start_addr_ctx1 = startAddr1[401:396]; 
assign MEMC66_burst_count_ctx1 = count1[468:462]; 
assign mAddr1[401:396] = MEMC66_addr_out_ctx1; 
assign mEn1[66:66] = MEMC66_mem_en_ctx1; 
assign mWEn1[66:66] = MEMC66_write_mem_en_ctx1; 
assign MEMC66_valid_ctx2 = valid2[66:66]; 
assign MEMC66_write_en_ctx2 = WEn2[66:66]; 
assign MEMC66_stride_ctx2 = stride2[66:66]; 
assign MEMC66_start_addr_ctx2 = startAddr2[401:396]; 
assign mAddr2[401:396] = MEMC66_addr_out_ctx2; 
assign MEMC66_burst_count_ctx2 = count2[468:462]; 
assign mEn2[66:66] = MEMC66_mem_en_ctx2; 
assign mWEn2[66:66] = MEMC66_write_mem_en_ctx2; 
wire [31:0] MEMOCMux67_inw1;
wire [31:0] MEMOCMux67_inw2;
wire [31:0] MEMOCMux67_inw3;
wire [31:0] MEMOCMux67_inw4;
wire [31:0] MEMOCMux67_inw5;
wire [31:0] MEMOCMux67_inw6;
wire [31:0] MEMOCMux67_inw7;
wire [31:0] MEMOCMux67_inw8;
wire [31:0] MEMOCMux67_inw9;
wire [31:0] MEMOCMux67_inw10;
wire [31:0] MEMOCMux67_outw1;
wire [3:0] MEMOCMux67_selw;
HA_10IM MEMOCMux67 (
.DataIn_1(MEMOCMux67_inw1),
.DataIn_2(MEMOCMux67_inw2),
.DataIn_3(MEMOCMux67_inw3),
.DataIn_4(MEMOCMux67_inw4),
.DataIn_5(MEMOCMux67_inw5),
.DataIn_6(MEMOCMux67_inw6),
.DataIn_7(MEMOCMux67_inw7),
.DataIn_8(MEMOCMux67_inw8),
.DataIn_9(MEMOCMux67_inw9),
.DataIn_10(MEMOCMux67_inw10),
.DataOut_1(MEMOCMux67_outw1),
.sel(MEMOCMux67_selw));
defparam MEMOCMux67.Mux_BW = 32;
assign MEMC67_data_from_Core = MEMOCMux67_outw1;
assign MEMOCMux67_inw1 = dataOutW[31:0]; 
assign MEMOCMux67_inw2 = dataOutW[63:32]; 
assign MEMOCMux67_inw3 = dataOutW[95:64]; 
assign MEMOCMux67_inw4 = dataOutW[127:96]; 
assign MEMOCMux67_inw5 = dataOutW[159:128]; 
assign MEMOCMux67_inw6 = dataOutW[191:160]; 
assign MEMOCMux67_inw7 = dataOutW[223:192]; 
assign MEMOCMux67_inw8 = dataOutW[255:224]; 
assign MEMOCMux67_inw9 = dataOutW[287:256]; 
assign MEMOCMux67_inw10 = globalDataIn[2175:2144]; 
assign MEMOCMux67_selw = mOutConfigW[271:268]; 
assign MEMC67_data_out_ctx2 = mDataFromMem[2175:2144]; 
assign mDataToMem[2175:2144] = MEMC67_data_in_ctx1; 
assign globalDataOut[2175:2144] = MEMC67_data_to_Core; 
assign MEMC67_valid_ctx1 = valid1[67:67]; 
assign MEMC67_write_en_ctx1 = WEn1[67:67]; 
assign MEMC67_stride_ctx1 = stride1[67:67]; 
assign MEMC67_start_addr_ctx1 = startAddr1[407:402]; 
assign MEMC67_burst_count_ctx1 = count1[475:469]; 
assign mAddr1[407:402] = MEMC67_addr_out_ctx1; 
assign mEn1[67:67] = MEMC67_mem_en_ctx1; 
assign mWEn1[67:67] = MEMC67_write_mem_en_ctx1; 
assign MEMC67_valid_ctx2 = valid2[67:67]; 
assign MEMC67_write_en_ctx2 = WEn2[67:67]; 
assign MEMC67_stride_ctx2 = stride2[67:67]; 
assign MEMC67_start_addr_ctx2 = startAddr2[407:402]; 
assign mAddr2[407:402] = MEMC67_addr_out_ctx2; 
assign MEMC67_burst_count_ctx2 = count2[475:469]; 
assign mEn2[67:67] = MEMC67_mem_en_ctx2; 
assign mWEn2[67:67] = MEMC67_write_mem_en_ctx2; 
wire [31:0] MEMOCMux68_inw1;
wire [31:0] MEMOCMux68_inw2;
wire [31:0] MEMOCMux68_inw3;
wire [31:0] MEMOCMux68_inw4;
wire [31:0] MEMOCMux68_inw5;
wire [31:0] MEMOCMux68_inw6;
wire [31:0] MEMOCMux68_inw7;
wire [31:0] MEMOCMux68_inw8;
wire [31:0] MEMOCMux68_inw9;
wire [31:0] MEMOCMux68_inw10;
wire [31:0] MEMOCMux68_outw1;
wire [3:0] MEMOCMux68_selw;
HA_10IM MEMOCMux68 (
.DataIn_1(MEMOCMux68_inw1),
.DataIn_2(MEMOCMux68_inw2),
.DataIn_3(MEMOCMux68_inw3),
.DataIn_4(MEMOCMux68_inw4),
.DataIn_5(MEMOCMux68_inw5),
.DataIn_6(MEMOCMux68_inw6),
.DataIn_7(MEMOCMux68_inw7),
.DataIn_8(MEMOCMux68_inw8),
.DataIn_9(MEMOCMux68_inw9),
.DataIn_10(MEMOCMux68_inw10),
.DataOut_1(MEMOCMux68_outw1),
.sel(MEMOCMux68_selw));
defparam MEMOCMux68.Mux_BW = 32;
assign MEMC68_data_from_Core = MEMOCMux68_outw1;
assign MEMOCMux68_inw1 = dataOutW[31:0]; 
assign MEMOCMux68_inw2 = dataOutW[63:32]; 
assign MEMOCMux68_inw3 = dataOutW[95:64]; 
assign MEMOCMux68_inw4 = dataOutW[127:96]; 
assign MEMOCMux68_inw5 = dataOutW[159:128]; 
assign MEMOCMux68_inw6 = dataOutW[191:160]; 
assign MEMOCMux68_inw7 = dataOutW[223:192]; 
assign MEMOCMux68_inw8 = dataOutW[255:224]; 
assign MEMOCMux68_inw9 = dataOutW[287:256]; 
assign MEMOCMux68_inw10 = globalDataIn[2207:2176]; 
assign MEMOCMux68_selw = mOutConfigW[275:272]; 
assign MEMC68_data_out_ctx2 = mDataFromMem[2207:2176]; 
assign mDataToMem[2207:2176] = MEMC68_data_in_ctx1; 
assign globalDataOut[2207:2176] = MEMC68_data_to_Core; 
assign MEMC68_valid_ctx1 = valid1[68:68]; 
assign MEMC68_write_en_ctx1 = WEn1[68:68]; 
assign MEMC68_stride_ctx1 = stride1[68:68]; 
assign MEMC68_start_addr_ctx1 = startAddr1[413:408]; 
assign MEMC68_burst_count_ctx1 = count1[482:476]; 
assign mAddr1[413:408] = MEMC68_addr_out_ctx1; 
assign mEn1[68:68] = MEMC68_mem_en_ctx1; 
assign mWEn1[68:68] = MEMC68_write_mem_en_ctx1; 
assign MEMC68_valid_ctx2 = valid2[68:68]; 
assign MEMC68_write_en_ctx2 = WEn2[68:68]; 
assign MEMC68_stride_ctx2 = stride2[68:68]; 
assign MEMC68_start_addr_ctx2 = startAddr2[413:408]; 
assign mAddr2[413:408] = MEMC68_addr_out_ctx2; 
assign MEMC68_burst_count_ctx2 = count2[482:476]; 
assign mEn2[68:68] = MEMC68_mem_en_ctx2; 
assign mWEn2[68:68] = MEMC68_write_mem_en_ctx2; 
wire [31:0] MEMOCMux69_inw1;
wire [31:0] MEMOCMux69_inw2;
wire [31:0] MEMOCMux69_inw3;
wire [31:0] MEMOCMux69_inw4;
wire [31:0] MEMOCMux69_inw5;
wire [31:0] MEMOCMux69_inw6;
wire [31:0] MEMOCMux69_inw7;
wire [31:0] MEMOCMux69_inw8;
wire [31:0] MEMOCMux69_inw9;
wire [31:0] MEMOCMux69_inw10;
wire [31:0] MEMOCMux69_outw1;
wire [3:0] MEMOCMux69_selw;
HA_10IM MEMOCMux69 (
.DataIn_1(MEMOCMux69_inw1),
.DataIn_2(MEMOCMux69_inw2),
.DataIn_3(MEMOCMux69_inw3),
.DataIn_4(MEMOCMux69_inw4),
.DataIn_5(MEMOCMux69_inw5),
.DataIn_6(MEMOCMux69_inw6),
.DataIn_7(MEMOCMux69_inw7),
.DataIn_8(MEMOCMux69_inw8),
.DataIn_9(MEMOCMux69_inw9),
.DataIn_10(MEMOCMux69_inw10),
.DataOut_1(MEMOCMux69_outw1),
.sel(MEMOCMux69_selw));
defparam MEMOCMux69.Mux_BW = 32;
assign MEMC69_data_from_Core = MEMOCMux69_outw1;
assign MEMOCMux69_inw1 = dataOutW[31:0]; 
assign MEMOCMux69_inw2 = dataOutW[63:32]; 
assign MEMOCMux69_inw3 = dataOutW[95:64]; 
assign MEMOCMux69_inw4 = dataOutW[127:96]; 
assign MEMOCMux69_inw5 = dataOutW[159:128]; 
assign MEMOCMux69_inw6 = dataOutW[191:160]; 
assign MEMOCMux69_inw7 = dataOutW[223:192]; 
assign MEMOCMux69_inw8 = dataOutW[255:224]; 
assign MEMOCMux69_inw9 = dataOutW[287:256]; 
assign MEMOCMux69_inw10 = globalDataIn[2239:2208]; 
assign MEMOCMux69_selw = mOutConfigW[279:276]; 
assign MEMC69_data_out_ctx2 = mDataFromMem[2239:2208]; 
assign mDataToMem[2239:2208] = MEMC69_data_in_ctx1; 
assign globalDataOut[2239:2208] = MEMC69_data_to_Core; 
assign MEMC69_valid_ctx1 = valid1[69:69]; 
assign MEMC69_write_en_ctx1 = WEn1[69:69]; 
assign MEMC69_stride_ctx1 = stride1[69:69]; 
assign MEMC69_start_addr_ctx1 = startAddr1[419:414]; 
assign MEMC69_burst_count_ctx1 = count1[489:483]; 
assign mAddr1[419:414] = MEMC69_addr_out_ctx1; 
assign mEn1[69:69] = MEMC69_mem_en_ctx1; 
assign mWEn1[69:69] = MEMC69_write_mem_en_ctx1; 
assign MEMC69_valid_ctx2 = valid2[69:69]; 
assign MEMC69_write_en_ctx2 = WEn2[69:69]; 
assign MEMC69_stride_ctx2 = stride2[69:69]; 
assign MEMC69_start_addr_ctx2 = startAddr2[419:414]; 
assign mAddr2[419:414] = MEMC69_addr_out_ctx2; 
assign MEMC69_burst_count_ctx2 = count2[489:483]; 
assign mEn2[69:69] = MEMC69_mem_en_ctx2; 
assign mWEn2[69:69] = MEMC69_write_mem_en_ctx2; 
wire [31:0] MEMOCMux70_inw1;
wire [31:0] MEMOCMux70_inw2;
wire [31:0] MEMOCMux70_inw3;
wire [31:0] MEMOCMux70_inw4;
wire [31:0] MEMOCMux70_inw5;
wire [31:0] MEMOCMux70_inw6;
wire [31:0] MEMOCMux70_inw7;
wire [31:0] MEMOCMux70_inw8;
wire [31:0] MEMOCMux70_inw9;
wire [31:0] MEMOCMux70_inw10;
wire [31:0] MEMOCMux70_outw1;
wire [3:0] MEMOCMux70_selw;
HA_10IM MEMOCMux70 (
.DataIn_1(MEMOCMux70_inw1),
.DataIn_2(MEMOCMux70_inw2),
.DataIn_3(MEMOCMux70_inw3),
.DataIn_4(MEMOCMux70_inw4),
.DataIn_5(MEMOCMux70_inw5),
.DataIn_6(MEMOCMux70_inw6),
.DataIn_7(MEMOCMux70_inw7),
.DataIn_8(MEMOCMux70_inw8),
.DataIn_9(MEMOCMux70_inw9),
.DataIn_10(MEMOCMux70_inw10),
.DataOut_1(MEMOCMux70_outw1),
.sel(MEMOCMux70_selw));
defparam MEMOCMux70.Mux_BW = 32;
assign MEMC70_data_from_Core = MEMOCMux70_outw1;
assign MEMOCMux70_inw1 = dataOutW[31:0]; 
assign MEMOCMux70_inw2 = dataOutW[63:32]; 
assign MEMOCMux70_inw3 = dataOutW[95:64]; 
assign MEMOCMux70_inw4 = dataOutW[127:96]; 
assign MEMOCMux70_inw5 = dataOutW[159:128]; 
assign MEMOCMux70_inw6 = dataOutW[191:160]; 
assign MEMOCMux70_inw7 = dataOutW[223:192]; 
assign MEMOCMux70_inw8 = dataOutW[255:224]; 
assign MEMOCMux70_inw9 = dataOutW[287:256]; 
assign MEMOCMux70_inw10 = globalDataIn[2271:2240]; 
assign MEMOCMux70_selw = mOutConfigW[283:280]; 
assign MEMC70_data_out_ctx2 = mDataFromMem[2271:2240]; 
assign mDataToMem[2271:2240] = MEMC70_data_in_ctx1; 
assign globalDataOut[2271:2240] = MEMC70_data_to_Core; 
assign MEMC70_valid_ctx1 = valid1[70:70]; 
assign MEMC70_write_en_ctx1 = WEn1[70:70]; 
assign MEMC70_stride_ctx1 = stride1[70:70]; 
assign MEMC70_start_addr_ctx1 = startAddr1[425:420]; 
assign MEMC70_burst_count_ctx1 = count1[496:490]; 
assign mAddr1[425:420] = MEMC70_addr_out_ctx1; 
assign mEn1[70:70] = MEMC70_mem_en_ctx1; 
assign mWEn1[70:70] = MEMC70_write_mem_en_ctx1; 
assign MEMC70_valid_ctx2 = valid2[70:70]; 
assign MEMC70_write_en_ctx2 = WEn2[70:70]; 
assign MEMC70_stride_ctx2 = stride2[70:70]; 
assign MEMC70_start_addr_ctx2 = startAddr2[425:420]; 
assign mAddr2[425:420] = MEMC70_addr_out_ctx2; 
assign MEMC70_burst_count_ctx2 = count2[496:490]; 
assign mEn2[70:70] = MEMC70_mem_en_ctx2; 
assign mWEn2[70:70] = MEMC70_write_mem_en_ctx2; 
wire [31:0] MEMOCMux71_inw1;
wire [31:0] MEMOCMux71_inw2;
wire [31:0] MEMOCMux71_inw3;
wire [31:0] MEMOCMux71_inw4;
wire [31:0] MEMOCMux71_inw5;
wire [31:0] MEMOCMux71_inw6;
wire [31:0] MEMOCMux71_inw7;
wire [31:0] MEMOCMux71_inw8;
wire [31:0] MEMOCMux71_inw9;
wire [31:0] MEMOCMux71_inw10;
wire [31:0] MEMOCMux71_outw1;
wire [3:0] MEMOCMux71_selw;
HA_10IM MEMOCMux71 (
.DataIn_1(MEMOCMux71_inw1),
.DataIn_2(MEMOCMux71_inw2),
.DataIn_3(MEMOCMux71_inw3),
.DataIn_4(MEMOCMux71_inw4),
.DataIn_5(MEMOCMux71_inw5),
.DataIn_6(MEMOCMux71_inw6),
.DataIn_7(MEMOCMux71_inw7),
.DataIn_8(MEMOCMux71_inw8),
.DataIn_9(MEMOCMux71_inw9),
.DataIn_10(MEMOCMux71_inw10),
.DataOut_1(MEMOCMux71_outw1),
.sel(MEMOCMux71_selw));
defparam MEMOCMux71.Mux_BW = 32;
assign MEMC71_data_from_Core = MEMOCMux71_outw1;
assign MEMOCMux71_inw1 = dataOutW[31:0]; 
assign MEMOCMux71_inw2 = dataOutW[63:32]; 
assign MEMOCMux71_inw3 = dataOutW[95:64]; 
assign MEMOCMux71_inw4 = dataOutW[127:96]; 
assign MEMOCMux71_inw5 = dataOutW[159:128]; 
assign MEMOCMux71_inw6 = dataOutW[191:160]; 
assign MEMOCMux71_inw7 = dataOutW[223:192]; 
assign MEMOCMux71_inw8 = dataOutW[255:224]; 
assign MEMOCMux71_inw9 = dataOutW[287:256]; 
assign MEMOCMux71_inw10 = globalDataIn[2303:2272]; 
assign MEMOCMux71_selw = mOutConfigW[287:284]; 
assign MEMC71_data_out_ctx2 = mDataFromMem[2303:2272]; 
assign mDataToMem[2303:2272] = MEMC71_data_in_ctx1; 
assign globalDataOut[2303:2272] = MEMC71_data_to_Core; 
assign MEMC71_valid_ctx1 = valid1[71:71]; 
assign MEMC71_write_en_ctx1 = WEn1[71:71]; 
assign MEMC71_stride_ctx1 = stride1[71:71]; 
assign MEMC71_start_addr_ctx1 = startAddr1[431:426]; 
assign MEMC71_burst_count_ctx1 = count1[503:497]; 
assign mAddr1[431:426] = MEMC71_addr_out_ctx1; 
assign mEn1[71:71] = MEMC71_mem_en_ctx1; 
assign mWEn1[71:71] = MEMC71_write_mem_en_ctx1; 
assign MEMC71_valid_ctx2 = valid2[71:71]; 
assign MEMC71_write_en_ctx2 = WEn2[71:71]; 
assign MEMC71_stride_ctx2 = stride2[71:71]; 
assign MEMC71_start_addr_ctx2 = startAddr2[431:426]; 
assign mAddr2[431:426] = MEMC71_addr_out_ctx2; 
assign MEMC71_burst_count_ctx2 = count2[503:497]; 
assign mEn2[71:71] = MEMC71_mem_en_ctx2; 
assign mWEn2[71:71] = MEMC71_write_mem_en_ctx2; 
wire [31:0] MEMOCMux72_inw1;
wire [31:0] MEMOCMux72_inw2;
wire [31:0] MEMOCMux72_inw3;
wire [31:0] MEMOCMux72_inw4;
wire [31:0] MEMOCMux72_inw5;
wire [31:0] MEMOCMux72_inw6;
wire [31:0] MEMOCMux72_inw7;
wire [31:0] MEMOCMux72_inw8;
wire [31:0] MEMOCMux72_inw9;
wire [31:0] MEMOCMux72_inw10;
wire [31:0] MEMOCMux72_outw1;
wire [3:0] MEMOCMux72_selw;
HA_10IM MEMOCMux72 (
.DataIn_1(MEMOCMux72_inw1),
.DataIn_2(MEMOCMux72_inw2),
.DataIn_3(MEMOCMux72_inw3),
.DataIn_4(MEMOCMux72_inw4),
.DataIn_5(MEMOCMux72_inw5),
.DataIn_6(MEMOCMux72_inw6),
.DataIn_7(MEMOCMux72_inw7),
.DataIn_8(MEMOCMux72_inw8),
.DataIn_9(MEMOCMux72_inw9),
.DataIn_10(MEMOCMux72_inw10),
.DataOut_1(MEMOCMux72_outw1),
.sel(MEMOCMux72_selw));
defparam MEMOCMux72.Mux_BW = 32;
assign MEMC72_data_from_Core = MEMOCMux72_outw1;
assign MEMOCMux72_inw1 = dataOutW[31:0]; 
assign MEMOCMux72_inw2 = dataOutW[63:32]; 
assign MEMOCMux72_inw3 = dataOutW[95:64]; 
assign MEMOCMux72_inw4 = dataOutW[127:96]; 
assign MEMOCMux72_inw5 = dataOutW[159:128]; 
assign MEMOCMux72_inw6 = dataOutW[191:160]; 
assign MEMOCMux72_inw7 = dataOutW[223:192]; 
assign MEMOCMux72_inw8 = dataOutW[255:224]; 
assign MEMOCMux72_inw9 = dataOutW[287:256]; 
assign MEMOCMux72_inw10 = globalDataIn[2335:2304]; 
assign MEMOCMux72_selw = mOutConfigW[291:288]; 
assign MEMC72_data_out_ctx2 = mDataFromMem[2335:2304]; 
assign mDataToMem[2335:2304] = MEMC72_data_in_ctx1; 
assign globalDataOut[2335:2304] = MEMC72_data_to_Core; 
assign MEMC72_valid_ctx1 = valid1[72:72]; 
assign MEMC72_write_en_ctx1 = WEn1[72:72]; 
assign MEMC72_stride_ctx1 = stride1[72:72]; 
assign MEMC72_start_addr_ctx1 = startAddr1[437:432]; 
assign MEMC72_burst_count_ctx1 = count1[510:504]; 
assign mAddr1[437:432] = MEMC72_addr_out_ctx1; 
assign mEn1[72:72] = MEMC72_mem_en_ctx1; 
assign mWEn1[72:72] = MEMC72_write_mem_en_ctx1; 
assign MEMC72_valid_ctx2 = valid2[72:72]; 
assign MEMC72_write_en_ctx2 = WEn2[72:72]; 
assign MEMC72_stride_ctx2 = stride2[72:72]; 
assign MEMC72_start_addr_ctx2 = startAddr2[437:432]; 
assign mAddr2[437:432] = MEMC72_addr_out_ctx2; 
assign MEMC72_burst_count_ctx2 = count2[510:504]; 
assign mEn2[72:72] = MEMC72_mem_en_ctx2; 
assign mWEn2[72:72] = MEMC72_write_mem_en_ctx2; 
wire [31:0] MEMOCMux73_inw1;
wire [31:0] MEMOCMux73_inw2;
wire [31:0] MEMOCMux73_inw3;
wire [31:0] MEMOCMux73_inw4;
wire [31:0] MEMOCMux73_inw5;
wire [31:0] MEMOCMux73_inw6;
wire [31:0] MEMOCMux73_inw7;
wire [31:0] MEMOCMux73_inw8;
wire [31:0] MEMOCMux73_inw9;
wire [31:0] MEMOCMux73_inw10;
wire [31:0] MEMOCMux73_outw1;
wire [3:0] MEMOCMux73_selw;
HA_10IM MEMOCMux73 (
.DataIn_1(MEMOCMux73_inw1),
.DataIn_2(MEMOCMux73_inw2),
.DataIn_3(MEMOCMux73_inw3),
.DataIn_4(MEMOCMux73_inw4),
.DataIn_5(MEMOCMux73_inw5),
.DataIn_6(MEMOCMux73_inw6),
.DataIn_7(MEMOCMux73_inw7),
.DataIn_8(MEMOCMux73_inw8),
.DataIn_9(MEMOCMux73_inw9),
.DataIn_10(MEMOCMux73_inw10),
.DataOut_1(MEMOCMux73_outw1),
.sel(MEMOCMux73_selw));
defparam MEMOCMux73.Mux_BW = 32;
assign MEMC73_data_from_Core = MEMOCMux73_outw1;
assign MEMOCMux73_inw1 = dataOutW[31:0]; 
assign MEMOCMux73_inw2 = dataOutW[63:32]; 
assign MEMOCMux73_inw3 = dataOutW[95:64]; 
assign MEMOCMux73_inw4 = dataOutW[127:96]; 
assign MEMOCMux73_inw5 = dataOutW[159:128]; 
assign MEMOCMux73_inw6 = dataOutW[191:160]; 
assign MEMOCMux73_inw7 = dataOutW[223:192]; 
assign MEMOCMux73_inw8 = dataOutW[255:224]; 
assign MEMOCMux73_inw9 = dataOutW[287:256]; 
assign MEMOCMux73_inw10 = globalDataIn[2367:2336]; 
assign MEMOCMux73_selw = mOutConfigW[295:292]; 
assign MEMC73_data_out_ctx2 = mDataFromMem[2367:2336]; 
assign mDataToMem[2367:2336] = MEMC73_data_in_ctx1; 
assign globalDataOut[2367:2336] = MEMC73_data_to_Core; 
assign MEMC73_valid_ctx1 = valid1[73:73]; 
assign MEMC73_write_en_ctx1 = WEn1[73:73]; 
assign MEMC73_stride_ctx1 = stride1[73:73]; 
assign MEMC73_start_addr_ctx1 = startAddr1[443:438]; 
assign MEMC73_burst_count_ctx1 = count1[517:511]; 
assign mAddr1[443:438] = MEMC73_addr_out_ctx1; 
assign mEn1[73:73] = MEMC73_mem_en_ctx1; 
assign mWEn1[73:73] = MEMC73_write_mem_en_ctx1; 
assign MEMC73_valid_ctx2 = valid2[73:73]; 
assign MEMC73_write_en_ctx2 = WEn2[73:73]; 
assign MEMC73_stride_ctx2 = stride2[73:73]; 
assign MEMC73_start_addr_ctx2 = startAddr2[443:438]; 
assign mAddr2[443:438] = MEMC73_addr_out_ctx2; 
assign MEMC73_burst_count_ctx2 = count2[517:511]; 
assign mEn2[73:73] = MEMC73_mem_en_ctx2; 
assign mWEn2[73:73] = MEMC73_write_mem_en_ctx2; 
wire [31:0] MEMOCMux74_inw1;
wire [31:0] MEMOCMux74_inw2;
wire [31:0] MEMOCMux74_inw3;
wire [31:0] MEMOCMux74_inw4;
wire [31:0] MEMOCMux74_inw5;
wire [31:0] MEMOCMux74_inw6;
wire [31:0] MEMOCMux74_inw7;
wire [31:0] MEMOCMux74_inw8;
wire [31:0] MEMOCMux74_inw9;
wire [31:0] MEMOCMux74_inw10;
wire [31:0] MEMOCMux74_outw1;
wire [3:0] MEMOCMux74_selw;
HA_10IM MEMOCMux74 (
.DataIn_1(MEMOCMux74_inw1),
.DataIn_2(MEMOCMux74_inw2),
.DataIn_3(MEMOCMux74_inw3),
.DataIn_4(MEMOCMux74_inw4),
.DataIn_5(MEMOCMux74_inw5),
.DataIn_6(MEMOCMux74_inw6),
.DataIn_7(MEMOCMux74_inw7),
.DataIn_8(MEMOCMux74_inw8),
.DataIn_9(MEMOCMux74_inw9),
.DataIn_10(MEMOCMux74_inw10),
.DataOut_1(MEMOCMux74_outw1),
.sel(MEMOCMux74_selw));
defparam MEMOCMux74.Mux_BW = 32;
assign MEMC74_data_from_Core = MEMOCMux74_outw1;
assign MEMOCMux74_inw1 = dataOutW[31:0]; 
assign MEMOCMux74_inw2 = dataOutW[63:32]; 
assign MEMOCMux74_inw3 = dataOutW[95:64]; 
assign MEMOCMux74_inw4 = dataOutW[127:96]; 
assign MEMOCMux74_inw5 = dataOutW[159:128]; 
assign MEMOCMux74_inw6 = dataOutW[191:160]; 
assign MEMOCMux74_inw7 = dataOutW[223:192]; 
assign MEMOCMux74_inw8 = dataOutW[255:224]; 
assign MEMOCMux74_inw9 = dataOutW[287:256]; 
assign MEMOCMux74_inw10 = globalDataIn[2399:2368]; 
assign MEMOCMux74_selw = mOutConfigW[299:296]; 
assign MEMC74_data_out_ctx2 = mDataFromMem[2399:2368]; 
assign mDataToMem[2399:2368] = MEMC74_data_in_ctx1; 
assign globalDataOut[2399:2368] = MEMC74_data_to_Core; 
assign MEMC74_valid_ctx1 = valid1[74:74]; 
assign MEMC74_write_en_ctx1 = WEn1[74:74]; 
assign MEMC74_stride_ctx1 = stride1[74:74]; 
assign MEMC74_start_addr_ctx1 = startAddr1[449:444]; 
assign MEMC74_burst_count_ctx1 = count1[524:518]; 
assign mAddr1[449:444] = MEMC74_addr_out_ctx1; 
assign mEn1[74:74] = MEMC74_mem_en_ctx1; 
assign mWEn1[74:74] = MEMC74_write_mem_en_ctx1; 
assign MEMC74_valid_ctx2 = valid2[74:74]; 
assign MEMC74_write_en_ctx2 = WEn2[74:74]; 
assign MEMC74_stride_ctx2 = stride2[74:74]; 
assign MEMC74_start_addr_ctx2 = startAddr2[449:444]; 
assign mAddr2[449:444] = MEMC74_addr_out_ctx2; 
assign MEMC74_burst_count_ctx2 = count2[524:518]; 
assign mEn2[74:74] = MEMC74_mem_en_ctx2; 
assign mWEn2[74:74] = MEMC74_write_mem_en_ctx2; 
wire [31:0] MEMOCMux75_inw1;
wire [31:0] MEMOCMux75_inw2;
wire [31:0] MEMOCMux75_inw3;
wire [31:0] MEMOCMux75_inw4;
wire [31:0] MEMOCMux75_inw5;
wire [31:0] MEMOCMux75_inw6;
wire [31:0] MEMOCMux75_inw7;
wire [31:0] MEMOCMux75_inw8;
wire [31:0] MEMOCMux75_inw9;
wire [31:0] MEMOCMux75_inw10;
wire [31:0] MEMOCMux75_outw1;
wire [3:0] MEMOCMux75_selw;
HA_10IM MEMOCMux75 (
.DataIn_1(MEMOCMux75_inw1),
.DataIn_2(MEMOCMux75_inw2),
.DataIn_3(MEMOCMux75_inw3),
.DataIn_4(MEMOCMux75_inw4),
.DataIn_5(MEMOCMux75_inw5),
.DataIn_6(MEMOCMux75_inw6),
.DataIn_7(MEMOCMux75_inw7),
.DataIn_8(MEMOCMux75_inw8),
.DataIn_9(MEMOCMux75_inw9),
.DataIn_10(MEMOCMux75_inw10),
.DataOut_1(MEMOCMux75_outw1),
.sel(MEMOCMux75_selw));
defparam MEMOCMux75.Mux_BW = 32;
assign MEMC75_data_from_Core = MEMOCMux75_outw1;
assign MEMOCMux75_inw1 = dataOutW[31:0]; 
assign MEMOCMux75_inw2 = dataOutW[63:32]; 
assign MEMOCMux75_inw3 = dataOutW[95:64]; 
assign MEMOCMux75_inw4 = dataOutW[127:96]; 
assign MEMOCMux75_inw5 = dataOutW[159:128]; 
assign MEMOCMux75_inw6 = dataOutW[191:160]; 
assign MEMOCMux75_inw7 = dataOutW[223:192]; 
assign MEMOCMux75_inw8 = dataOutW[255:224]; 
assign MEMOCMux75_inw9 = dataOutW[287:256]; 
assign MEMOCMux75_inw10 = globalDataIn[2431:2400]; 
assign MEMOCMux75_selw = mOutConfigW[303:300]; 
assign MEMC75_data_out_ctx2 = mDataFromMem[2431:2400]; 
assign mDataToMem[2431:2400] = MEMC75_data_in_ctx1; 
assign globalDataOut[2431:2400] = MEMC75_data_to_Core; 
assign MEMC75_valid_ctx1 = valid1[75:75]; 
assign MEMC75_write_en_ctx1 = WEn1[75:75]; 
assign MEMC75_stride_ctx1 = stride1[75:75]; 
assign MEMC75_start_addr_ctx1 = startAddr1[455:450]; 
assign MEMC75_burst_count_ctx1 = count1[531:525]; 
assign mAddr1[455:450] = MEMC75_addr_out_ctx1; 
assign mEn1[75:75] = MEMC75_mem_en_ctx1; 
assign mWEn1[75:75] = MEMC75_write_mem_en_ctx1; 
assign MEMC75_valid_ctx2 = valid2[75:75]; 
assign MEMC75_write_en_ctx2 = WEn2[75:75]; 
assign MEMC75_stride_ctx2 = stride2[75:75]; 
assign MEMC75_start_addr_ctx2 = startAddr2[455:450]; 
assign mAddr2[455:450] = MEMC75_addr_out_ctx2; 
assign MEMC75_burst_count_ctx2 = count2[531:525]; 
assign mEn2[75:75] = MEMC75_mem_en_ctx2; 
assign mWEn2[75:75] = MEMC75_write_mem_en_ctx2; 
wire [31:0] MEMOCMux76_inw1;
wire [31:0] MEMOCMux76_inw2;
wire [31:0] MEMOCMux76_inw3;
wire [31:0] MEMOCMux76_inw4;
wire [31:0] MEMOCMux76_inw5;
wire [31:0] MEMOCMux76_inw6;
wire [31:0] MEMOCMux76_inw7;
wire [31:0] MEMOCMux76_inw8;
wire [31:0] MEMOCMux76_inw9;
wire [31:0] MEMOCMux76_inw10;
wire [31:0] MEMOCMux76_outw1;
wire [3:0] MEMOCMux76_selw;
HA_10IM MEMOCMux76 (
.DataIn_1(MEMOCMux76_inw1),
.DataIn_2(MEMOCMux76_inw2),
.DataIn_3(MEMOCMux76_inw3),
.DataIn_4(MEMOCMux76_inw4),
.DataIn_5(MEMOCMux76_inw5),
.DataIn_6(MEMOCMux76_inw6),
.DataIn_7(MEMOCMux76_inw7),
.DataIn_8(MEMOCMux76_inw8),
.DataIn_9(MEMOCMux76_inw9),
.DataIn_10(MEMOCMux76_inw10),
.DataOut_1(MEMOCMux76_outw1),
.sel(MEMOCMux76_selw));
defparam MEMOCMux76.Mux_BW = 32;
assign MEMC76_data_from_Core = MEMOCMux76_outw1;
assign MEMOCMux76_inw1 = dataOutW[31:0]; 
assign MEMOCMux76_inw2 = dataOutW[63:32]; 
assign MEMOCMux76_inw3 = dataOutW[95:64]; 
assign MEMOCMux76_inw4 = dataOutW[127:96]; 
assign MEMOCMux76_inw5 = dataOutW[159:128]; 
assign MEMOCMux76_inw6 = dataOutW[191:160]; 
assign MEMOCMux76_inw7 = dataOutW[223:192]; 
assign MEMOCMux76_inw8 = dataOutW[255:224]; 
assign MEMOCMux76_inw9 = dataOutW[287:256]; 
assign MEMOCMux76_inw10 = globalDataIn[2463:2432]; 
assign MEMOCMux76_selw = mOutConfigW[307:304]; 
assign MEMC76_data_out_ctx2 = mDataFromMem[2463:2432]; 
assign mDataToMem[2463:2432] = MEMC76_data_in_ctx1; 
assign globalDataOut[2463:2432] = MEMC76_data_to_Core; 
assign MEMC76_valid_ctx1 = valid1[76:76]; 
assign MEMC76_write_en_ctx1 = WEn1[76:76]; 
assign MEMC76_stride_ctx1 = stride1[76:76]; 
assign MEMC76_start_addr_ctx1 = startAddr1[461:456]; 
assign MEMC76_burst_count_ctx1 = count1[538:532]; 
assign mAddr1[461:456] = MEMC76_addr_out_ctx1; 
assign mEn1[76:76] = MEMC76_mem_en_ctx1; 
assign mWEn1[76:76] = MEMC76_write_mem_en_ctx1; 
assign MEMC76_valid_ctx2 = valid2[76:76]; 
assign MEMC76_write_en_ctx2 = WEn2[76:76]; 
assign MEMC76_stride_ctx2 = stride2[76:76]; 
assign MEMC76_start_addr_ctx2 = startAddr2[461:456]; 
assign mAddr2[461:456] = MEMC76_addr_out_ctx2; 
assign MEMC76_burst_count_ctx2 = count2[538:532]; 
assign mEn2[76:76] = MEMC76_mem_en_ctx2; 
assign mWEn2[76:76] = MEMC76_write_mem_en_ctx2; 
wire [31:0] MEMOCMux77_inw1;
wire [31:0] MEMOCMux77_inw2;
wire [31:0] MEMOCMux77_inw3;
wire [31:0] MEMOCMux77_inw4;
wire [31:0] MEMOCMux77_inw5;
wire [31:0] MEMOCMux77_inw6;
wire [31:0] MEMOCMux77_inw7;
wire [31:0] MEMOCMux77_inw8;
wire [31:0] MEMOCMux77_inw9;
wire [31:0] MEMOCMux77_inw10;
wire [31:0] MEMOCMux77_outw1;
wire [3:0] MEMOCMux77_selw;
HA_10IM MEMOCMux77 (
.DataIn_1(MEMOCMux77_inw1),
.DataIn_2(MEMOCMux77_inw2),
.DataIn_3(MEMOCMux77_inw3),
.DataIn_4(MEMOCMux77_inw4),
.DataIn_5(MEMOCMux77_inw5),
.DataIn_6(MEMOCMux77_inw6),
.DataIn_7(MEMOCMux77_inw7),
.DataIn_8(MEMOCMux77_inw8),
.DataIn_9(MEMOCMux77_inw9),
.DataIn_10(MEMOCMux77_inw10),
.DataOut_1(MEMOCMux77_outw1),
.sel(MEMOCMux77_selw));
defparam MEMOCMux77.Mux_BW = 32;
assign MEMC77_data_from_Core = MEMOCMux77_outw1;
assign MEMOCMux77_inw1 = dataOutW[31:0]; 
assign MEMOCMux77_inw2 = dataOutW[63:32]; 
assign MEMOCMux77_inw3 = dataOutW[95:64]; 
assign MEMOCMux77_inw4 = dataOutW[127:96]; 
assign MEMOCMux77_inw5 = dataOutW[159:128]; 
assign MEMOCMux77_inw6 = dataOutW[191:160]; 
assign MEMOCMux77_inw7 = dataOutW[223:192]; 
assign MEMOCMux77_inw8 = dataOutW[255:224]; 
assign MEMOCMux77_inw9 = dataOutW[287:256]; 
assign MEMOCMux77_inw10 = globalDataIn[2495:2464]; 
assign MEMOCMux77_selw = mOutConfigW[311:308]; 
assign MEMC77_data_out_ctx2 = mDataFromMem[2495:2464]; 
assign mDataToMem[2495:2464] = MEMC77_data_in_ctx1; 
assign globalDataOut[2495:2464] = MEMC77_data_to_Core; 
assign MEMC77_valid_ctx1 = valid1[77:77]; 
assign MEMC77_write_en_ctx1 = WEn1[77:77]; 
assign MEMC77_stride_ctx1 = stride1[77:77]; 
assign MEMC77_start_addr_ctx1 = startAddr1[467:462]; 
assign MEMC77_burst_count_ctx1 = count1[545:539]; 
assign mAddr1[467:462] = MEMC77_addr_out_ctx1; 
assign mEn1[77:77] = MEMC77_mem_en_ctx1; 
assign mWEn1[77:77] = MEMC77_write_mem_en_ctx1; 
assign MEMC77_valid_ctx2 = valid2[77:77]; 
assign MEMC77_write_en_ctx2 = WEn2[77:77]; 
assign MEMC77_stride_ctx2 = stride2[77:77]; 
assign MEMC77_start_addr_ctx2 = startAddr2[467:462]; 
assign mAddr2[467:462] = MEMC77_addr_out_ctx2; 
assign MEMC77_burst_count_ctx2 = count2[545:539]; 
assign mEn2[77:77] = MEMC77_mem_en_ctx2; 
assign mWEn2[77:77] = MEMC77_write_mem_en_ctx2; 
wire [31:0] MEMOCMux78_inw1;
wire [31:0] MEMOCMux78_inw2;
wire [31:0] MEMOCMux78_inw3;
wire [31:0] MEMOCMux78_inw4;
wire [31:0] MEMOCMux78_inw5;
wire [31:0] MEMOCMux78_inw6;
wire [31:0] MEMOCMux78_inw7;
wire [31:0] MEMOCMux78_inw8;
wire [31:0] MEMOCMux78_inw9;
wire [31:0] MEMOCMux78_inw10;
wire [31:0] MEMOCMux78_outw1;
wire [3:0] MEMOCMux78_selw;
HA_10IM MEMOCMux78 (
.DataIn_1(MEMOCMux78_inw1),
.DataIn_2(MEMOCMux78_inw2),
.DataIn_3(MEMOCMux78_inw3),
.DataIn_4(MEMOCMux78_inw4),
.DataIn_5(MEMOCMux78_inw5),
.DataIn_6(MEMOCMux78_inw6),
.DataIn_7(MEMOCMux78_inw7),
.DataIn_8(MEMOCMux78_inw8),
.DataIn_9(MEMOCMux78_inw9),
.DataIn_10(MEMOCMux78_inw10),
.DataOut_1(MEMOCMux78_outw1),
.sel(MEMOCMux78_selw));
defparam MEMOCMux78.Mux_BW = 32;
assign MEMC78_data_from_Core = MEMOCMux78_outw1;
assign MEMOCMux78_inw1 = dataOutW[31:0]; 
assign MEMOCMux78_inw2 = dataOutW[63:32]; 
assign MEMOCMux78_inw3 = dataOutW[95:64]; 
assign MEMOCMux78_inw4 = dataOutW[127:96]; 
assign MEMOCMux78_inw5 = dataOutW[159:128]; 
assign MEMOCMux78_inw6 = dataOutW[191:160]; 
assign MEMOCMux78_inw7 = dataOutW[223:192]; 
assign MEMOCMux78_inw8 = dataOutW[255:224]; 
assign MEMOCMux78_inw9 = dataOutW[287:256]; 
assign MEMOCMux78_inw10 = globalDataIn[2527:2496]; 
assign MEMOCMux78_selw = mOutConfigW[315:312]; 
assign MEMC78_data_out_ctx2 = mDataFromMem[2527:2496]; 
assign mDataToMem[2527:2496] = MEMC78_data_in_ctx1; 
assign globalDataOut[2527:2496] = MEMC78_data_to_Core; 
assign MEMC78_valid_ctx1 = valid1[78:78]; 
assign MEMC78_write_en_ctx1 = WEn1[78:78]; 
assign MEMC78_stride_ctx1 = stride1[78:78]; 
assign MEMC78_start_addr_ctx1 = startAddr1[473:468]; 
assign MEMC78_burst_count_ctx1 = count1[552:546]; 
assign mAddr1[473:468] = MEMC78_addr_out_ctx1; 
assign mEn1[78:78] = MEMC78_mem_en_ctx1; 
assign mWEn1[78:78] = MEMC78_write_mem_en_ctx1; 
assign MEMC78_valid_ctx2 = valid2[78:78]; 
assign MEMC78_write_en_ctx2 = WEn2[78:78]; 
assign MEMC78_stride_ctx2 = stride2[78:78]; 
assign MEMC78_start_addr_ctx2 = startAddr2[473:468]; 
assign mAddr2[473:468] = MEMC78_addr_out_ctx2; 
assign MEMC78_burst_count_ctx2 = count2[552:546]; 
assign mEn2[78:78] = MEMC78_mem_en_ctx2; 
assign mWEn2[78:78] = MEMC78_write_mem_en_ctx2; 
wire [31:0] MEMOCMux79_inw1;
wire [31:0] MEMOCMux79_inw2;
wire [31:0] MEMOCMux79_inw3;
wire [31:0] MEMOCMux79_inw4;
wire [31:0] MEMOCMux79_inw5;
wire [31:0] MEMOCMux79_inw6;
wire [31:0] MEMOCMux79_inw7;
wire [31:0] MEMOCMux79_inw8;
wire [31:0] MEMOCMux79_inw9;
wire [31:0] MEMOCMux79_inw10;
wire [31:0] MEMOCMux79_outw1;
wire [3:0] MEMOCMux79_selw;
HA_10IM MEMOCMux79 (
.DataIn_1(MEMOCMux79_inw1),
.DataIn_2(MEMOCMux79_inw2),
.DataIn_3(MEMOCMux79_inw3),
.DataIn_4(MEMOCMux79_inw4),
.DataIn_5(MEMOCMux79_inw5),
.DataIn_6(MEMOCMux79_inw6),
.DataIn_7(MEMOCMux79_inw7),
.DataIn_8(MEMOCMux79_inw8),
.DataIn_9(MEMOCMux79_inw9),
.DataIn_10(MEMOCMux79_inw10),
.DataOut_1(MEMOCMux79_outw1),
.sel(MEMOCMux79_selw));
defparam MEMOCMux79.Mux_BW = 32;
assign MEMC79_data_from_Core = MEMOCMux79_outw1;
assign MEMOCMux79_inw1 = dataOutW[31:0]; 
assign MEMOCMux79_inw2 = dataOutW[63:32]; 
assign MEMOCMux79_inw3 = dataOutW[95:64]; 
assign MEMOCMux79_inw4 = dataOutW[127:96]; 
assign MEMOCMux79_inw5 = dataOutW[159:128]; 
assign MEMOCMux79_inw6 = dataOutW[191:160]; 
assign MEMOCMux79_inw7 = dataOutW[223:192]; 
assign MEMOCMux79_inw8 = dataOutW[255:224]; 
assign MEMOCMux79_inw9 = dataOutW[287:256]; 
assign MEMOCMux79_inw10 = globalDataIn[2559:2528]; 
assign MEMOCMux79_selw = mOutConfigW[319:316]; 
assign MEMC79_data_out_ctx2 = mDataFromMem[2559:2528]; 
assign mDataToMem[2559:2528] = MEMC79_data_in_ctx1; 
assign globalDataOut[2559:2528] = MEMC79_data_to_Core; 
assign MEMC79_valid_ctx1 = valid1[79:79]; 
assign MEMC79_write_en_ctx1 = WEn1[79:79]; 
assign MEMC79_stride_ctx1 = stride1[79:79]; 
assign MEMC79_start_addr_ctx1 = startAddr1[479:474]; 
assign MEMC79_burst_count_ctx1 = count1[559:553]; 
assign mAddr1[479:474] = MEMC79_addr_out_ctx1; 
assign mEn1[79:79] = MEMC79_mem_en_ctx1; 
assign mWEn1[79:79] = MEMC79_write_mem_en_ctx1; 
assign MEMC79_valid_ctx2 = valid2[79:79]; 
assign MEMC79_write_en_ctx2 = WEn2[79:79]; 
assign MEMC79_stride_ctx2 = stride2[79:79]; 
assign MEMC79_start_addr_ctx2 = startAddr2[479:474]; 
assign mAddr2[479:474] = MEMC79_addr_out_ctx2; 
assign MEMC79_burst_count_ctx2 = count2[559:553]; 
assign mEn2[79:79] = MEMC79_mem_en_ctx2; 
assign mWEn2[79:79] = MEMC79_write_mem_en_ctx2; 
wire [31:0] MEMOCMux80_inw1;
wire [31:0] MEMOCMux80_inw2;
wire [31:0] MEMOCMux80_inw3;
wire [31:0] MEMOCMux80_inw4;
wire [31:0] MEMOCMux80_inw5;
wire [31:0] MEMOCMux80_inw6;
wire [31:0] MEMOCMux80_inw7;
wire [31:0] MEMOCMux80_inw8;
wire [31:0] MEMOCMux80_inw9;
wire [31:0] MEMOCMux80_inw10;
wire [31:0] MEMOCMux80_outw1;
wire [3:0] MEMOCMux80_selw;
HA_10IM MEMOCMux80 (
.DataIn_1(MEMOCMux80_inw1),
.DataIn_2(MEMOCMux80_inw2),
.DataIn_3(MEMOCMux80_inw3),
.DataIn_4(MEMOCMux80_inw4),
.DataIn_5(MEMOCMux80_inw5),
.DataIn_6(MEMOCMux80_inw6),
.DataIn_7(MEMOCMux80_inw7),
.DataIn_8(MEMOCMux80_inw8),
.DataIn_9(MEMOCMux80_inw9),
.DataIn_10(MEMOCMux80_inw10),
.DataOut_1(MEMOCMux80_outw1),
.sel(MEMOCMux80_selw));
defparam MEMOCMux80.Mux_BW = 32;
assign MEMC80_data_from_Core = MEMOCMux80_outw1;
assign MEMOCMux80_inw1 = dataOutW[31:0]; 
assign MEMOCMux80_inw2 = dataOutW[63:32]; 
assign MEMOCMux80_inw3 = dataOutW[95:64]; 
assign MEMOCMux80_inw4 = dataOutW[127:96]; 
assign MEMOCMux80_inw5 = dataOutW[159:128]; 
assign MEMOCMux80_inw6 = dataOutW[191:160]; 
assign MEMOCMux80_inw7 = dataOutW[223:192]; 
assign MEMOCMux80_inw8 = dataOutW[255:224]; 
assign MEMOCMux80_inw9 = dataOutW[287:256]; 
assign MEMOCMux80_inw10 = globalDataIn[2591:2560]; 
assign MEMOCMux80_selw = mOutConfigW[323:320]; 
assign MEMC80_data_out_ctx2 = mDataFromMem[2591:2560]; 
assign mDataToMem[2591:2560] = MEMC80_data_in_ctx1; 
assign globalDataOut[2591:2560] = MEMC80_data_to_Core; 
assign MEMC80_valid_ctx1 = valid1[80:80]; 
assign MEMC80_write_en_ctx1 = WEn1[80:80]; 
assign MEMC80_stride_ctx1 = stride1[80:80]; 
assign MEMC80_start_addr_ctx1 = startAddr1[485:480]; 
assign MEMC80_burst_count_ctx1 = count1[566:560]; 
assign mAddr1[485:480] = MEMC80_addr_out_ctx1; 
assign mEn1[80:80] = MEMC80_mem_en_ctx1; 
assign mWEn1[80:80] = MEMC80_write_mem_en_ctx1; 
assign MEMC80_valid_ctx2 = valid2[80:80]; 
assign MEMC80_write_en_ctx2 = WEn2[80:80]; 
assign MEMC80_stride_ctx2 = stride2[80:80]; 
assign MEMC80_start_addr_ctx2 = startAddr2[485:480]; 
assign mAddr2[485:480] = MEMC80_addr_out_ctx2; 
assign MEMC80_burst_count_ctx2 = count2[566:560]; 
assign mEn2[80:80] = MEMC80_mem_en_ctx2; 
assign mWEn2[80:80] = MEMC80_write_mem_en_ctx2; 
wire [31:0] MEMOCMux81_inw1;
wire [31:0] MEMOCMux81_inw2;
wire [31:0] MEMOCMux81_inw3;
wire [31:0] MEMOCMux81_inw4;
wire [31:0] MEMOCMux81_inw5;
wire [31:0] MEMOCMux81_inw6;
wire [31:0] MEMOCMux81_inw7;
wire [31:0] MEMOCMux81_inw8;
wire [31:0] MEMOCMux81_inw9;
wire [31:0] MEMOCMux81_inw10;
wire [31:0] MEMOCMux81_outw1;
wire [3:0] MEMOCMux81_selw;
HA_10IM MEMOCMux81 (
.DataIn_1(MEMOCMux81_inw1),
.DataIn_2(MEMOCMux81_inw2),
.DataIn_3(MEMOCMux81_inw3),
.DataIn_4(MEMOCMux81_inw4),
.DataIn_5(MEMOCMux81_inw5),
.DataIn_6(MEMOCMux81_inw6),
.DataIn_7(MEMOCMux81_inw7),
.DataIn_8(MEMOCMux81_inw8),
.DataIn_9(MEMOCMux81_inw9),
.DataIn_10(MEMOCMux81_inw10),
.DataOut_1(MEMOCMux81_outw1),
.sel(MEMOCMux81_selw));
defparam MEMOCMux81.Mux_BW = 32;
assign MEMC81_data_from_Core = MEMOCMux81_outw1;
assign MEMOCMux81_inw1 = dataOutW[31:0]; 
assign MEMOCMux81_inw2 = dataOutW[63:32]; 
assign MEMOCMux81_inw3 = dataOutW[95:64]; 
assign MEMOCMux81_inw4 = dataOutW[127:96]; 
assign MEMOCMux81_inw5 = dataOutW[159:128]; 
assign MEMOCMux81_inw6 = dataOutW[191:160]; 
assign MEMOCMux81_inw7 = dataOutW[223:192]; 
assign MEMOCMux81_inw8 = dataOutW[255:224]; 
assign MEMOCMux81_inw9 = dataOutW[287:256]; 
assign MEMOCMux81_inw10 = globalDataIn[2623:2592]; 
assign MEMOCMux81_selw = mOutConfigW[327:324]; 
assign MEMC81_data_out_ctx2 = mDataFromMem[2623:2592]; 
assign mDataToMem[2623:2592] = MEMC81_data_in_ctx1; 
assign globalDataOut[2623:2592] = MEMC81_data_to_Core; 
assign MEMC81_valid_ctx1 = valid1[81:81]; 
assign MEMC81_write_en_ctx1 = WEn1[81:81]; 
assign MEMC81_stride_ctx1 = stride1[81:81]; 
assign MEMC81_start_addr_ctx1 = startAddr1[491:486]; 
assign MEMC81_burst_count_ctx1 = count1[573:567]; 
assign mAddr1[491:486] = MEMC81_addr_out_ctx1; 
assign mEn1[81:81] = MEMC81_mem_en_ctx1; 
assign mWEn1[81:81] = MEMC81_write_mem_en_ctx1; 
assign MEMC81_valid_ctx2 = valid2[81:81]; 
assign MEMC81_write_en_ctx2 = WEn2[81:81]; 
assign MEMC81_stride_ctx2 = stride2[81:81]; 
assign MEMC81_start_addr_ctx2 = startAddr2[491:486]; 
assign mAddr2[491:486] = MEMC81_addr_out_ctx2; 
assign MEMC81_burst_count_ctx2 = count2[573:567]; 
assign mEn2[81:81] = MEMC81_mem_en_ctx2; 
assign mWEn2[81:81] = MEMC81_write_mem_en_ctx2; 
wire [31:0] MEMOCMux82_inw1;
wire [31:0] MEMOCMux82_inw2;
wire [31:0] MEMOCMux82_inw3;
wire [31:0] MEMOCMux82_inw4;
wire [31:0] MEMOCMux82_inw5;
wire [31:0] MEMOCMux82_inw6;
wire [31:0] MEMOCMux82_inw7;
wire [31:0] MEMOCMux82_inw8;
wire [31:0] MEMOCMux82_inw9;
wire [31:0] MEMOCMux82_inw10;
wire [31:0] MEMOCMux82_outw1;
wire [3:0] MEMOCMux82_selw;
HA_10IM MEMOCMux82 (
.DataIn_1(MEMOCMux82_inw1),
.DataIn_2(MEMOCMux82_inw2),
.DataIn_3(MEMOCMux82_inw3),
.DataIn_4(MEMOCMux82_inw4),
.DataIn_5(MEMOCMux82_inw5),
.DataIn_6(MEMOCMux82_inw6),
.DataIn_7(MEMOCMux82_inw7),
.DataIn_8(MEMOCMux82_inw8),
.DataIn_9(MEMOCMux82_inw9),
.DataIn_10(MEMOCMux82_inw10),
.DataOut_1(MEMOCMux82_outw1),
.sel(MEMOCMux82_selw));
defparam MEMOCMux82.Mux_BW = 32;
assign MEMC82_data_from_Core = MEMOCMux82_outw1;
assign MEMOCMux82_inw1 = dataOutW[31:0]; 
assign MEMOCMux82_inw2 = dataOutW[63:32]; 
assign MEMOCMux82_inw3 = dataOutW[95:64]; 
assign MEMOCMux82_inw4 = dataOutW[127:96]; 
assign MEMOCMux82_inw5 = dataOutW[159:128]; 
assign MEMOCMux82_inw6 = dataOutW[191:160]; 
assign MEMOCMux82_inw7 = dataOutW[223:192]; 
assign MEMOCMux82_inw8 = dataOutW[255:224]; 
assign MEMOCMux82_inw9 = dataOutW[287:256]; 
assign MEMOCMux82_inw10 = globalDataIn[2655:2624]; 
assign MEMOCMux82_selw = mOutConfigW[331:328]; 
assign MEMC82_data_out_ctx2 = mDataFromMem[2655:2624]; 
assign mDataToMem[2655:2624] = MEMC82_data_in_ctx1; 
assign globalDataOut[2655:2624] = MEMC82_data_to_Core; 
assign MEMC82_valid_ctx1 = valid1[82:82]; 
assign MEMC82_write_en_ctx1 = WEn1[82:82]; 
assign MEMC82_stride_ctx1 = stride1[82:82]; 
assign MEMC82_start_addr_ctx1 = startAddr1[497:492]; 
assign MEMC82_burst_count_ctx1 = count1[580:574]; 
assign mAddr1[497:492] = MEMC82_addr_out_ctx1; 
assign mEn1[82:82] = MEMC82_mem_en_ctx1; 
assign mWEn1[82:82] = MEMC82_write_mem_en_ctx1; 
assign MEMC82_valid_ctx2 = valid2[82:82]; 
assign MEMC82_write_en_ctx2 = WEn2[82:82]; 
assign MEMC82_stride_ctx2 = stride2[82:82]; 
assign MEMC82_start_addr_ctx2 = startAddr2[497:492]; 
assign mAddr2[497:492] = MEMC82_addr_out_ctx2; 
assign MEMC82_burst_count_ctx2 = count2[580:574]; 
assign mEn2[82:82] = MEMC82_mem_en_ctx2; 
assign mWEn2[82:82] = MEMC82_write_mem_en_ctx2; 
wire [31:0] MEMOCMux83_inw1;
wire [31:0] MEMOCMux83_inw2;
wire [31:0] MEMOCMux83_inw3;
wire [31:0] MEMOCMux83_inw4;
wire [31:0] MEMOCMux83_inw5;
wire [31:0] MEMOCMux83_inw6;
wire [31:0] MEMOCMux83_inw7;
wire [31:0] MEMOCMux83_inw8;
wire [31:0] MEMOCMux83_inw9;
wire [31:0] MEMOCMux83_inw10;
wire [31:0] MEMOCMux83_outw1;
wire [3:0] MEMOCMux83_selw;
HA_10IM MEMOCMux83 (
.DataIn_1(MEMOCMux83_inw1),
.DataIn_2(MEMOCMux83_inw2),
.DataIn_3(MEMOCMux83_inw3),
.DataIn_4(MEMOCMux83_inw4),
.DataIn_5(MEMOCMux83_inw5),
.DataIn_6(MEMOCMux83_inw6),
.DataIn_7(MEMOCMux83_inw7),
.DataIn_8(MEMOCMux83_inw8),
.DataIn_9(MEMOCMux83_inw9),
.DataIn_10(MEMOCMux83_inw10),
.DataOut_1(MEMOCMux83_outw1),
.sel(MEMOCMux83_selw));
defparam MEMOCMux83.Mux_BW = 32;
assign MEMC83_data_from_Core = MEMOCMux83_outw1;
assign MEMOCMux83_inw1 = dataOutW[31:0]; 
assign MEMOCMux83_inw2 = dataOutW[63:32]; 
assign MEMOCMux83_inw3 = dataOutW[95:64]; 
assign MEMOCMux83_inw4 = dataOutW[127:96]; 
assign MEMOCMux83_inw5 = dataOutW[159:128]; 
assign MEMOCMux83_inw6 = dataOutW[191:160]; 
assign MEMOCMux83_inw7 = dataOutW[223:192]; 
assign MEMOCMux83_inw8 = dataOutW[255:224]; 
assign MEMOCMux83_inw9 = dataOutW[287:256]; 
assign MEMOCMux83_inw10 = globalDataIn[2687:2656]; 
assign MEMOCMux83_selw = mOutConfigW[335:332]; 
assign MEMC83_data_out_ctx2 = mDataFromMem[2687:2656]; 
assign mDataToMem[2687:2656] = MEMC83_data_in_ctx1; 
assign globalDataOut[2687:2656] = MEMC83_data_to_Core; 
assign MEMC83_valid_ctx1 = valid1[83:83]; 
assign MEMC83_write_en_ctx1 = WEn1[83:83]; 
assign MEMC83_stride_ctx1 = stride1[83:83]; 
assign MEMC83_start_addr_ctx1 = startAddr1[503:498]; 
assign MEMC83_burst_count_ctx1 = count1[587:581]; 
assign mAddr1[503:498] = MEMC83_addr_out_ctx1; 
assign mEn1[83:83] = MEMC83_mem_en_ctx1; 
assign mWEn1[83:83] = MEMC83_write_mem_en_ctx1; 
assign MEMC83_valid_ctx2 = valid2[83:83]; 
assign MEMC83_write_en_ctx2 = WEn2[83:83]; 
assign MEMC83_stride_ctx2 = stride2[83:83]; 
assign MEMC83_start_addr_ctx2 = startAddr2[503:498]; 
assign mAddr2[503:498] = MEMC83_addr_out_ctx2; 
assign MEMC83_burst_count_ctx2 = count2[587:581]; 
assign mEn2[83:83] = MEMC83_mem_en_ctx2; 
assign mWEn2[83:83] = MEMC83_write_mem_en_ctx2; 
wire [31:0] MEMOCMux84_inw1;
wire [31:0] MEMOCMux84_inw2;
wire [31:0] MEMOCMux84_inw3;
wire [31:0] MEMOCMux84_inw4;
wire [31:0] MEMOCMux84_inw5;
wire [31:0] MEMOCMux84_inw6;
wire [31:0] MEMOCMux84_inw7;
wire [31:0] MEMOCMux84_inw8;
wire [31:0] MEMOCMux84_inw9;
wire [31:0] MEMOCMux84_inw10;
wire [31:0] MEMOCMux84_outw1;
wire [3:0] MEMOCMux84_selw;
HA_10IM MEMOCMux84 (
.DataIn_1(MEMOCMux84_inw1),
.DataIn_2(MEMOCMux84_inw2),
.DataIn_3(MEMOCMux84_inw3),
.DataIn_4(MEMOCMux84_inw4),
.DataIn_5(MEMOCMux84_inw5),
.DataIn_6(MEMOCMux84_inw6),
.DataIn_7(MEMOCMux84_inw7),
.DataIn_8(MEMOCMux84_inw8),
.DataIn_9(MEMOCMux84_inw9),
.DataIn_10(MEMOCMux84_inw10),
.DataOut_1(MEMOCMux84_outw1),
.sel(MEMOCMux84_selw));
defparam MEMOCMux84.Mux_BW = 32;
assign MEMC84_data_from_Core = MEMOCMux84_outw1;
assign MEMOCMux84_inw1 = dataOutW[31:0]; 
assign MEMOCMux84_inw2 = dataOutW[63:32]; 
assign MEMOCMux84_inw3 = dataOutW[95:64]; 
assign MEMOCMux84_inw4 = dataOutW[127:96]; 
assign MEMOCMux84_inw5 = dataOutW[159:128]; 
assign MEMOCMux84_inw6 = dataOutW[191:160]; 
assign MEMOCMux84_inw7 = dataOutW[223:192]; 
assign MEMOCMux84_inw8 = dataOutW[255:224]; 
assign MEMOCMux84_inw9 = dataOutW[287:256]; 
assign MEMOCMux84_inw10 = globalDataIn[2719:2688]; 
assign MEMOCMux84_selw = mOutConfigW[339:336]; 
assign MEMC84_data_out_ctx2 = mDataFromMem[2719:2688]; 
assign mDataToMem[2719:2688] = MEMC84_data_in_ctx1; 
assign globalDataOut[2719:2688] = MEMC84_data_to_Core; 
assign MEMC84_valid_ctx1 = valid1[84:84]; 
assign MEMC84_write_en_ctx1 = WEn1[84:84]; 
assign MEMC84_stride_ctx1 = stride1[84:84]; 
assign MEMC84_start_addr_ctx1 = startAddr1[509:504]; 
assign MEMC84_burst_count_ctx1 = count1[594:588]; 
assign mAddr1[509:504] = MEMC84_addr_out_ctx1; 
assign mEn1[84:84] = MEMC84_mem_en_ctx1; 
assign mWEn1[84:84] = MEMC84_write_mem_en_ctx1; 
assign MEMC84_valid_ctx2 = valid2[84:84]; 
assign MEMC84_write_en_ctx2 = WEn2[84:84]; 
assign MEMC84_stride_ctx2 = stride2[84:84]; 
assign MEMC84_start_addr_ctx2 = startAddr2[509:504]; 
assign mAddr2[509:504] = MEMC84_addr_out_ctx2; 
assign MEMC84_burst_count_ctx2 = count2[594:588]; 
assign mEn2[84:84] = MEMC84_mem_en_ctx2; 
assign mWEn2[84:84] = MEMC84_write_mem_en_ctx2; 
wire [31:0] MEMOCMux85_inw1;
wire [31:0] MEMOCMux85_inw2;
wire [31:0] MEMOCMux85_inw3;
wire [31:0] MEMOCMux85_inw4;
wire [31:0] MEMOCMux85_inw5;
wire [31:0] MEMOCMux85_inw6;
wire [31:0] MEMOCMux85_inw7;
wire [31:0] MEMOCMux85_inw8;
wire [31:0] MEMOCMux85_inw9;
wire [31:0] MEMOCMux85_inw10;
wire [31:0] MEMOCMux85_outw1;
wire [3:0] MEMOCMux85_selw;
HA_10IM MEMOCMux85 (
.DataIn_1(MEMOCMux85_inw1),
.DataIn_2(MEMOCMux85_inw2),
.DataIn_3(MEMOCMux85_inw3),
.DataIn_4(MEMOCMux85_inw4),
.DataIn_5(MEMOCMux85_inw5),
.DataIn_6(MEMOCMux85_inw6),
.DataIn_7(MEMOCMux85_inw7),
.DataIn_8(MEMOCMux85_inw8),
.DataIn_9(MEMOCMux85_inw9),
.DataIn_10(MEMOCMux85_inw10),
.DataOut_1(MEMOCMux85_outw1),
.sel(MEMOCMux85_selw));
defparam MEMOCMux85.Mux_BW = 32;
assign MEMC85_data_from_Core = MEMOCMux85_outw1;
assign MEMOCMux85_inw1 = dataOutW[31:0]; 
assign MEMOCMux85_inw2 = dataOutW[63:32]; 
assign MEMOCMux85_inw3 = dataOutW[95:64]; 
assign MEMOCMux85_inw4 = dataOutW[127:96]; 
assign MEMOCMux85_inw5 = dataOutW[159:128]; 
assign MEMOCMux85_inw6 = dataOutW[191:160]; 
assign MEMOCMux85_inw7 = dataOutW[223:192]; 
assign MEMOCMux85_inw8 = dataOutW[255:224]; 
assign MEMOCMux85_inw9 = dataOutW[287:256]; 
assign MEMOCMux85_inw10 = globalDataIn[2751:2720]; 
assign MEMOCMux85_selw = mOutConfigW[343:340]; 
assign MEMC85_data_out_ctx2 = mDataFromMem[2751:2720]; 
assign mDataToMem[2751:2720] = MEMC85_data_in_ctx1; 
assign globalDataOut[2751:2720] = MEMC85_data_to_Core; 
assign MEMC85_valid_ctx1 = valid1[85:85]; 
assign MEMC85_write_en_ctx1 = WEn1[85:85]; 
assign MEMC85_stride_ctx1 = stride1[85:85]; 
assign MEMC85_start_addr_ctx1 = startAddr1[515:510]; 
assign MEMC85_burst_count_ctx1 = count1[601:595]; 
assign mAddr1[515:510] = MEMC85_addr_out_ctx1; 
assign mEn1[85:85] = MEMC85_mem_en_ctx1; 
assign mWEn1[85:85] = MEMC85_write_mem_en_ctx1; 
assign MEMC85_valid_ctx2 = valid2[85:85]; 
assign MEMC85_write_en_ctx2 = WEn2[85:85]; 
assign MEMC85_stride_ctx2 = stride2[85:85]; 
assign MEMC85_start_addr_ctx2 = startAddr2[515:510]; 
assign mAddr2[515:510] = MEMC85_addr_out_ctx2; 
assign MEMC85_burst_count_ctx2 = count2[601:595]; 
assign mEn2[85:85] = MEMC85_mem_en_ctx2; 
assign mWEn2[85:85] = MEMC85_write_mem_en_ctx2; 
wire [31:0] MEMOCMux86_inw1;
wire [31:0] MEMOCMux86_inw2;
wire [31:0] MEMOCMux86_inw3;
wire [31:0] MEMOCMux86_inw4;
wire [31:0] MEMOCMux86_inw5;
wire [31:0] MEMOCMux86_inw6;
wire [31:0] MEMOCMux86_inw7;
wire [31:0] MEMOCMux86_inw8;
wire [31:0] MEMOCMux86_inw9;
wire [31:0] MEMOCMux86_inw10;
wire [31:0] MEMOCMux86_outw1;
wire [3:0] MEMOCMux86_selw;
HA_10IM MEMOCMux86 (
.DataIn_1(MEMOCMux86_inw1),
.DataIn_2(MEMOCMux86_inw2),
.DataIn_3(MEMOCMux86_inw3),
.DataIn_4(MEMOCMux86_inw4),
.DataIn_5(MEMOCMux86_inw5),
.DataIn_6(MEMOCMux86_inw6),
.DataIn_7(MEMOCMux86_inw7),
.DataIn_8(MEMOCMux86_inw8),
.DataIn_9(MEMOCMux86_inw9),
.DataIn_10(MEMOCMux86_inw10),
.DataOut_1(MEMOCMux86_outw1),
.sel(MEMOCMux86_selw));
defparam MEMOCMux86.Mux_BW = 32;
assign MEMC86_data_from_Core = MEMOCMux86_outw1;
assign MEMOCMux86_inw1 = dataOutW[31:0]; 
assign MEMOCMux86_inw2 = dataOutW[63:32]; 
assign MEMOCMux86_inw3 = dataOutW[95:64]; 
assign MEMOCMux86_inw4 = dataOutW[127:96]; 
assign MEMOCMux86_inw5 = dataOutW[159:128]; 
assign MEMOCMux86_inw6 = dataOutW[191:160]; 
assign MEMOCMux86_inw7 = dataOutW[223:192]; 
assign MEMOCMux86_inw8 = dataOutW[255:224]; 
assign MEMOCMux86_inw9 = dataOutW[287:256]; 
assign MEMOCMux86_inw10 = globalDataIn[2783:2752]; 
assign MEMOCMux86_selw = mOutConfigW[347:344]; 
assign MEMC86_data_out_ctx2 = mDataFromMem[2783:2752]; 
assign mDataToMem[2783:2752] = MEMC86_data_in_ctx1; 
assign globalDataOut[2783:2752] = MEMC86_data_to_Core; 
assign MEMC86_valid_ctx1 = valid1[86:86]; 
assign MEMC86_write_en_ctx1 = WEn1[86:86]; 
assign MEMC86_stride_ctx1 = stride1[86:86]; 
assign MEMC86_start_addr_ctx1 = startAddr1[521:516]; 
assign MEMC86_burst_count_ctx1 = count1[608:602]; 
assign mAddr1[521:516] = MEMC86_addr_out_ctx1; 
assign mEn1[86:86] = MEMC86_mem_en_ctx1; 
assign mWEn1[86:86] = MEMC86_write_mem_en_ctx1; 
assign MEMC86_valid_ctx2 = valid2[86:86]; 
assign MEMC86_write_en_ctx2 = WEn2[86:86]; 
assign MEMC86_stride_ctx2 = stride2[86:86]; 
assign MEMC86_start_addr_ctx2 = startAddr2[521:516]; 
assign mAddr2[521:516] = MEMC86_addr_out_ctx2; 
assign MEMC86_burst_count_ctx2 = count2[608:602]; 
assign mEn2[86:86] = MEMC86_mem_en_ctx2; 
assign mWEn2[86:86] = MEMC86_write_mem_en_ctx2; 
wire [31:0] MEMOCMux87_inw1;
wire [31:0] MEMOCMux87_inw2;
wire [31:0] MEMOCMux87_inw3;
wire [31:0] MEMOCMux87_inw4;
wire [31:0] MEMOCMux87_inw5;
wire [31:0] MEMOCMux87_inw6;
wire [31:0] MEMOCMux87_inw7;
wire [31:0] MEMOCMux87_inw8;
wire [31:0] MEMOCMux87_inw9;
wire [31:0] MEMOCMux87_inw10;
wire [31:0] MEMOCMux87_outw1;
wire [3:0] MEMOCMux87_selw;
HA_10IM MEMOCMux87 (
.DataIn_1(MEMOCMux87_inw1),
.DataIn_2(MEMOCMux87_inw2),
.DataIn_3(MEMOCMux87_inw3),
.DataIn_4(MEMOCMux87_inw4),
.DataIn_5(MEMOCMux87_inw5),
.DataIn_6(MEMOCMux87_inw6),
.DataIn_7(MEMOCMux87_inw7),
.DataIn_8(MEMOCMux87_inw8),
.DataIn_9(MEMOCMux87_inw9),
.DataIn_10(MEMOCMux87_inw10),
.DataOut_1(MEMOCMux87_outw1),
.sel(MEMOCMux87_selw));
defparam MEMOCMux87.Mux_BW = 32;
assign MEMC87_data_from_Core = MEMOCMux87_outw1;
assign MEMOCMux87_inw1 = dataOutW[31:0]; 
assign MEMOCMux87_inw2 = dataOutW[63:32]; 
assign MEMOCMux87_inw3 = dataOutW[95:64]; 
assign MEMOCMux87_inw4 = dataOutW[127:96]; 
assign MEMOCMux87_inw5 = dataOutW[159:128]; 
assign MEMOCMux87_inw6 = dataOutW[191:160]; 
assign MEMOCMux87_inw7 = dataOutW[223:192]; 
assign MEMOCMux87_inw8 = dataOutW[255:224]; 
assign MEMOCMux87_inw9 = dataOutW[287:256]; 
assign MEMOCMux87_inw10 = globalDataIn[2815:2784]; 
assign MEMOCMux87_selw = mOutConfigW[351:348]; 
assign MEMC87_data_out_ctx2 = mDataFromMem[2815:2784]; 
assign mDataToMem[2815:2784] = MEMC87_data_in_ctx1; 
assign globalDataOut[2815:2784] = MEMC87_data_to_Core; 
assign MEMC87_valid_ctx1 = valid1[87:87]; 
assign MEMC87_write_en_ctx1 = WEn1[87:87]; 
assign MEMC87_stride_ctx1 = stride1[87:87]; 
assign MEMC87_start_addr_ctx1 = startAddr1[527:522]; 
assign MEMC87_burst_count_ctx1 = count1[615:609]; 
assign mAddr1[527:522] = MEMC87_addr_out_ctx1; 
assign mEn1[87:87] = MEMC87_mem_en_ctx1; 
assign mWEn1[87:87] = MEMC87_write_mem_en_ctx1; 
assign MEMC87_valid_ctx2 = valid2[87:87]; 
assign MEMC87_write_en_ctx2 = WEn2[87:87]; 
assign MEMC87_stride_ctx2 = stride2[87:87]; 
assign MEMC87_start_addr_ctx2 = startAddr2[527:522]; 
assign mAddr2[527:522] = MEMC87_addr_out_ctx2; 
assign MEMC87_burst_count_ctx2 = count2[615:609]; 
assign mEn2[87:87] = MEMC87_mem_en_ctx2; 
assign mWEn2[87:87] = MEMC87_write_mem_en_ctx2; 
wire [31:0] MEMOCMux88_inw1;
wire [31:0] MEMOCMux88_inw2;
wire [31:0] MEMOCMux88_inw3;
wire [31:0] MEMOCMux88_inw4;
wire [31:0] MEMOCMux88_inw5;
wire [31:0] MEMOCMux88_inw6;
wire [31:0] MEMOCMux88_inw7;
wire [31:0] MEMOCMux88_inw8;
wire [31:0] MEMOCMux88_inw9;
wire [31:0] MEMOCMux88_inw10;
wire [31:0] MEMOCMux88_outw1;
wire [3:0] MEMOCMux88_selw;
HA_10IM MEMOCMux88 (
.DataIn_1(MEMOCMux88_inw1),
.DataIn_2(MEMOCMux88_inw2),
.DataIn_3(MEMOCMux88_inw3),
.DataIn_4(MEMOCMux88_inw4),
.DataIn_5(MEMOCMux88_inw5),
.DataIn_6(MEMOCMux88_inw6),
.DataIn_7(MEMOCMux88_inw7),
.DataIn_8(MEMOCMux88_inw8),
.DataIn_9(MEMOCMux88_inw9),
.DataIn_10(MEMOCMux88_inw10),
.DataOut_1(MEMOCMux88_outw1),
.sel(MEMOCMux88_selw));
defparam MEMOCMux88.Mux_BW = 32;
assign MEMC88_data_from_Core = MEMOCMux88_outw1;
assign MEMOCMux88_inw1 = dataOutW[31:0]; 
assign MEMOCMux88_inw2 = dataOutW[63:32]; 
assign MEMOCMux88_inw3 = dataOutW[95:64]; 
assign MEMOCMux88_inw4 = dataOutW[127:96]; 
assign MEMOCMux88_inw5 = dataOutW[159:128]; 
assign MEMOCMux88_inw6 = dataOutW[191:160]; 
assign MEMOCMux88_inw7 = dataOutW[223:192]; 
assign MEMOCMux88_inw8 = dataOutW[255:224]; 
assign MEMOCMux88_inw9 = dataOutW[287:256]; 
assign MEMOCMux88_inw10 = globalDataIn[2847:2816]; 
assign MEMOCMux88_selw = mOutConfigW[355:352]; 
assign MEMC88_data_out_ctx2 = mDataFromMem[2847:2816]; 
assign mDataToMem[2847:2816] = MEMC88_data_in_ctx1; 
assign globalDataOut[2847:2816] = MEMC88_data_to_Core; 
assign MEMC88_valid_ctx1 = valid1[88:88]; 
assign MEMC88_write_en_ctx1 = WEn1[88:88]; 
assign MEMC88_stride_ctx1 = stride1[88:88]; 
assign MEMC88_start_addr_ctx1 = startAddr1[533:528]; 
assign MEMC88_burst_count_ctx1 = count1[622:616]; 
assign mAddr1[533:528] = MEMC88_addr_out_ctx1; 
assign mEn1[88:88] = MEMC88_mem_en_ctx1; 
assign mWEn1[88:88] = MEMC88_write_mem_en_ctx1; 
assign MEMC88_valid_ctx2 = valid2[88:88]; 
assign MEMC88_write_en_ctx2 = WEn2[88:88]; 
assign MEMC88_stride_ctx2 = stride2[88:88]; 
assign MEMC88_start_addr_ctx2 = startAddr2[533:528]; 
assign mAddr2[533:528] = MEMC88_addr_out_ctx2; 
assign MEMC88_burst_count_ctx2 = count2[622:616]; 
assign mEn2[88:88] = MEMC88_mem_en_ctx2; 
assign mWEn2[88:88] = MEMC88_write_mem_en_ctx2; 
wire [31:0] MEMOCMux89_inw1;
wire [31:0] MEMOCMux89_inw2;
wire [31:0] MEMOCMux89_inw3;
wire [31:0] MEMOCMux89_inw4;
wire [31:0] MEMOCMux89_inw5;
wire [31:0] MEMOCMux89_inw6;
wire [31:0] MEMOCMux89_inw7;
wire [31:0] MEMOCMux89_inw8;
wire [31:0] MEMOCMux89_inw9;
wire [31:0] MEMOCMux89_inw10;
wire [31:0] MEMOCMux89_outw1;
wire [3:0] MEMOCMux89_selw;
HA_10IM MEMOCMux89 (
.DataIn_1(MEMOCMux89_inw1),
.DataIn_2(MEMOCMux89_inw2),
.DataIn_3(MEMOCMux89_inw3),
.DataIn_4(MEMOCMux89_inw4),
.DataIn_5(MEMOCMux89_inw5),
.DataIn_6(MEMOCMux89_inw6),
.DataIn_7(MEMOCMux89_inw7),
.DataIn_8(MEMOCMux89_inw8),
.DataIn_9(MEMOCMux89_inw9),
.DataIn_10(MEMOCMux89_inw10),
.DataOut_1(MEMOCMux89_outw1),
.sel(MEMOCMux89_selw));
defparam MEMOCMux89.Mux_BW = 32;
assign MEMC89_data_from_Core = MEMOCMux89_outw1;
assign MEMOCMux89_inw1 = dataOutW[31:0]; 
assign MEMOCMux89_inw2 = dataOutW[63:32]; 
assign MEMOCMux89_inw3 = dataOutW[95:64]; 
assign MEMOCMux89_inw4 = dataOutW[127:96]; 
assign MEMOCMux89_inw5 = dataOutW[159:128]; 
assign MEMOCMux89_inw6 = dataOutW[191:160]; 
assign MEMOCMux89_inw7 = dataOutW[223:192]; 
assign MEMOCMux89_inw8 = dataOutW[255:224]; 
assign MEMOCMux89_inw9 = dataOutW[287:256]; 
assign MEMOCMux89_inw10 = globalDataIn[2879:2848]; 
assign MEMOCMux89_selw = mOutConfigW[359:356]; 
assign MEMC89_data_out_ctx2 = mDataFromMem[2879:2848]; 
assign mDataToMem[2879:2848] = MEMC89_data_in_ctx1; 
assign globalDataOut[2879:2848] = MEMC89_data_to_Core; 
assign MEMC89_valid_ctx1 = valid1[89:89]; 
assign MEMC89_write_en_ctx1 = WEn1[89:89]; 
assign MEMC89_stride_ctx1 = stride1[89:89]; 
assign MEMC89_start_addr_ctx1 = startAddr1[539:534]; 
assign MEMC89_burst_count_ctx1 = count1[629:623]; 
assign mAddr1[539:534] = MEMC89_addr_out_ctx1; 
assign mEn1[89:89] = MEMC89_mem_en_ctx1; 
assign mWEn1[89:89] = MEMC89_write_mem_en_ctx1; 
assign MEMC89_valid_ctx2 = valid2[89:89]; 
assign MEMC89_write_en_ctx2 = WEn2[89:89]; 
assign MEMC89_stride_ctx2 = stride2[89:89]; 
assign MEMC89_start_addr_ctx2 = startAddr2[539:534]; 
assign mAddr2[539:534] = MEMC89_addr_out_ctx2; 
assign MEMC89_burst_count_ctx2 = count2[629:623]; 
assign mEn2[89:89] = MEMC89_mem_en_ctx2; 
assign mWEn2[89:89] = MEMC89_write_mem_en_ctx2; 
wire [31:0] MEMOCMux90_inw1;
wire [31:0] MEMOCMux90_inw2;
wire [31:0] MEMOCMux90_inw3;
wire [31:0] MEMOCMux90_inw4;
wire [31:0] MEMOCMux90_inw5;
wire [31:0] MEMOCMux90_inw6;
wire [31:0] MEMOCMux90_inw7;
wire [31:0] MEMOCMux90_inw8;
wire [31:0] MEMOCMux90_inw9;
wire [31:0] MEMOCMux90_inw10;
wire [31:0] MEMOCMux90_outw1;
wire [3:0] MEMOCMux90_selw;
HA_10IM MEMOCMux90 (
.DataIn_1(MEMOCMux90_inw1),
.DataIn_2(MEMOCMux90_inw2),
.DataIn_3(MEMOCMux90_inw3),
.DataIn_4(MEMOCMux90_inw4),
.DataIn_5(MEMOCMux90_inw5),
.DataIn_6(MEMOCMux90_inw6),
.DataIn_7(MEMOCMux90_inw7),
.DataIn_8(MEMOCMux90_inw8),
.DataIn_9(MEMOCMux90_inw9),
.DataIn_10(MEMOCMux90_inw10),
.DataOut_1(MEMOCMux90_outw1),
.sel(MEMOCMux90_selw));
defparam MEMOCMux90.Mux_BW = 32;
assign MEMC90_data_from_Core = MEMOCMux90_outw1;
assign MEMOCMux90_inw1 = dataOutW[31:0]; 
assign MEMOCMux90_inw2 = dataOutW[63:32]; 
assign MEMOCMux90_inw3 = dataOutW[95:64]; 
assign MEMOCMux90_inw4 = dataOutW[127:96]; 
assign MEMOCMux90_inw5 = dataOutW[159:128]; 
assign MEMOCMux90_inw6 = dataOutW[191:160]; 
assign MEMOCMux90_inw7 = dataOutW[223:192]; 
assign MEMOCMux90_inw8 = dataOutW[255:224]; 
assign MEMOCMux90_inw9 = dataOutW[287:256]; 
assign MEMOCMux90_inw10 = globalDataIn[2911:2880]; 
assign MEMOCMux90_selw = mOutConfigW[363:360]; 
assign MEMC90_data_out_ctx2 = mDataFromMem[2911:2880]; 
assign mDataToMem[2911:2880] = MEMC90_data_in_ctx1; 
assign globalDataOut[2911:2880] = MEMC90_data_to_Core; 
assign MEMC90_valid_ctx1 = valid1[90:90]; 
assign MEMC90_write_en_ctx1 = WEn1[90:90]; 
assign MEMC90_stride_ctx1 = stride1[90:90]; 
assign MEMC90_start_addr_ctx1 = startAddr1[545:540]; 
assign MEMC90_burst_count_ctx1 = count1[636:630]; 
assign mAddr1[545:540] = MEMC90_addr_out_ctx1; 
assign mEn1[90:90] = MEMC90_mem_en_ctx1; 
assign mWEn1[90:90] = MEMC90_write_mem_en_ctx1; 
assign MEMC90_valid_ctx2 = valid2[90:90]; 
assign MEMC90_write_en_ctx2 = WEn2[90:90]; 
assign MEMC90_stride_ctx2 = stride2[90:90]; 
assign MEMC90_start_addr_ctx2 = startAddr2[545:540]; 
assign mAddr2[545:540] = MEMC90_addr_out_ctx2; 
assign MEMC90_burst_count_ctx2 = count2[636:630]; 
assign mEn2[90:90] = MEMC90_mem_en_ctx2; 
assign mWEn2[90:90] = MEMC90_write_mem_en_ctx2; 
wire [31:0] MEMOCMux91_inw1;
wire [31:0] MEMOCMux91_inw2;
wire [31:0] MEMOCMux91_inw3;
wire [31:0] MEMOCMux91_inw4;
wire [31:0] MEMOCMux91_inw5;
wire [31:0] MEMOCMux91_inw6;
wire [31:0] MEMOCMux91_inw7;
wire [31:0] MEMOCMux91_inw8;
wire [31:0] MEMOCMux91_inw9;
wire [31:0] MEMOCMux91_inw10;
wire [31:0] MEMOCMux91_outw1;
wire [3:0] MEMOCMux91_selw;
HA_10IM MEMOCMux91 (
.DataIn_1(MEMOCMux91_inw1),
.DataIn_2(MEMOCMux91_inw2),
.DataIn_3(MEMOCMux91_inw3),
.DataIn_4(MEMOCMux91_inw4),
.DataIn_5(MEMOCMux91_inw5),
.DataIn_6(MEMOCMux91_inw6),
.DataIn_7(MEMOCMux91_inw7),
.DataIn_8(MEMOCMux91_inw8),
.DataIn_9(MEMOCMux91_inw9),
.DataIn_10(MEMOCMux91_inw10),
.DataOut_1(MEMOCMux91_outw1),
.sel(MEMOCMux91_selw));
defparam MEMOCMux91.Mux_BW = 32;
assign MEMC91_data_from_Core = MEMOCMux91_outw1;
assign MEMOCMux91_inw1 = dataOutW[31:0]; 
assign MEMOCMux91_inw2 = dataOutW[63:32]; 
assign MEMOCMux91_inw3 = dataOutW[95:64]; 
assign MEMOCMux91_inw4 = dataOutW[127:96]; 
assign MEMOCMux91_inw5 = dataOutW[159:128]; 
assign MEMOCMux91_inw6 = dataOutW[191:160]; 
assign MEMOCMux91_inw7 = dataOutW[223:192]; 
assign MEMOCMux91_inw8 = dataOutW[255:224]; 
assign MEMOCMux91_inw9 = dataOutW[287:256]; 
assign MEMOCMux91_inw10 = globalDataIn[2943:2912]; 
assign MEMOCMux91_selw = mOutConfigW[367:364]; 
assign MEMC91_data_out_ctx2 = mDataFromMem[2943:2912]; 
assign mDataToMem[2943:2912] = MEMC91_data_in_ctx1; 
assign globalDataOut[2943:2912] = MEMC91_data_to_Core; 
assign MEMC91_valid_ctx1 = valid1[91:91]; 
assign MEMC91_write_en_ctx1 = WEn1[91:91]; 
assign MEMC91_stride_ctx1 = stride1[91:91]; 
assign MEMC91_start_addr_ctx1 = startAddr1[551:546]; 
assign MEMC91_burst_count_ctx1 = count1[643:637]; 
assign mAddr1[551:546] = MEMC91_addr_out_ctx1; 
assign mEn1[91:91] = MEMC91_mem_en_ctx1; 
assign mWEn1[91:91] = MEMC91_write_mem_en_ctx1; 
assign MEMC91_valid_ctx2 = valid2[91:91]; 
assign MEMC91_write_en_ctx2 = WEn2[91:91]; 
assign MEMC91_stride_ctx2 = stride2[91:91]; 
assign MEMC91_start_addr_ctx2 = startAddr2[551:546]; 
assign mAddr2[551:546] = MEMC91_addr_out_ctx2; 
assign MEMC91_burst_count_ctx2 = count2[643:637]; 
assign mEn2[91:91] = MEMC91_mem_en_ctx2; 
assign mWEn2[91:91] = MEMC91_write_mem_en_ctx2; 
wire [31:0] MEMOCMux92_inw1;
wire [31:0] MEMOCMux92_inw2;
wire [31:0] MEMOCMux92_inw3;
wire [31:0] MEMOCMux92_inw4;
wire [31:0] MEMOCMux92_inw5;
wire [31:0] MEMOCMux92_inw6;
wire [31:0] MEMOCMux92_inw7;
wire [31:0] MEMOCMux92_inw8;
wire [31:0] MEMOCMux92_inw9;
wire [31:0] MEMOCMux92_inw10;
wire [31:0] MEMOCMux92_outw1;
wire [3:0] MEMOCMux92_selw;
HA_10IM MEMOCMux92 (
.DataIn_1(MEMOCMux92_inw1),
.DataIn_2(MEMOCMux92_inw2),
.DataIn_3(MEMOCMux92_inw3),
.DataIn_4(MEMOCMux92_inw4),
.DataIn_5(MEMOCMux92_inw5),
.DataIn_6(MEMOCMux92_inw6),
.DataIn_7(MEMOCMux92_inw7),
.DataIn_8(MEMOCMux92_inw8),
.DataIn_9(MEMOCMux92_inw9),
.DataIn_10(MEMOCMux92_inw10),
.DataOut_1(MEMOCMux92_outw1),
.sel(MEMOCMux92_selw));
defparam MEMOCMux92.Mux_BW = 32;
assign MEMC92_data_from_Core = MEMOCMux92_outw1;
assign MEMOCMux92_inw1 = dataOutW[31:0]; 
assign MEMOCMux92_inw2 = dataOutW[63:32]; 
assign MEMOCMux92_inw3 = dataOutW[95:64]; 
assign MEMOCMux92_inw4 = dataOutW[127:96]; 
assign MEMOCMux92_inw5 = dataOutW[159:128]; 
assign MEMOCMux92_inw6 = dataOutW[191:160]; 
assign MEMOCMux92_inw7 = dataOutW[223:192]; 
assign MEMOCMux92_inw8 = dataOutW[255:224]; 
assign MEMOCMux92_inw9 = dataOutW[287:256]; 
assign MEMOCMux92_inw10 = globalDataIn[2975:2944]; 
assign MEMOCMux92_selw = mOutConfigW[371:368]; 
assign MEMC92_data_out_ctx2 = mDataFromMem[2975:2944]; 
assign mDataToMem[2975:2944] = MEMC92_data_in_ctx1; 
assign globalDataOut[2975:2944] = MEMC92_data_to_Core; 
assign MEMC92_valid_ctx1 = valid1[92:92]; 
assign MEMC92_write_en_ctx1 = WEn1[92:92]; 
assign MEMC92_stride_ctx1 = stride1[92:92]; 
assign MEMC92_start_addr_ctx1 = startAddr1[557:552]; 
assign MEMC92_burst_count_ctx1 = count1[650:644]; 
assign mAddr1[557:552] = MEMC92_addr_out_ctx1; 
assign mEn1[92:92] = MEMC92_mem_en_ctx1; 
assign mWEn1[92:92] = MEMC92_write_mem_en_ctx1; 
assign MEMC92_valid_ctx2 = valid2[92:92]; 
assign MEMC92_write_en_ctx2 = WEn2[92:92]; 
assign MEMC92_stride_ctx2 = stride2[92:92]; 
assign MEMC92_start_addr_ctx2 = startAddr2[557:552]; 
assign mAddr2[557:552] = MEMC92_addr_out_ctx2; 
assign MEMC92_burst_count_ctx2 = count2[650:644]; 
assign mEn2[92:92] = MEMC92_mem_en_ctx2; 
assign mWEn2[92:92] = MEMC92_write_mem_en_ctx2; 
wire [31:0] MEMOCMux93_inw1;
wire [31:0] MEMOCMux93_inw2;
wire [31:0] MEMOCMux93_inw3;
wire [31:0] MEMOCMux93_inw4;
wire [31:0] MEMOCMux93_inw5;
wire [31:0] MEMOCMux93_inw6;
wire [31:0] MEMOCMux93_inw7;
wire [31:0] MEMOCMux93_inw8;
wire [31:0] MEMOCMux93_inw9;
wire [31:0] MEMOCMux93_inw10;
wire [31:0] MEMOCMux93_outw1;
wire [3:0] MEMOCMux93_selw;
HA_10IM MEMOCMux93 (
.DataIn_1(MEMOCMux93_inw1),
.DataIn_2(MEMOCMux93_inw2),
.DataIn_3(MEMOCMux93_inw3),
.DataIn_4(MEMOCMux93_inw4),
.DataIn_5(MEMOCMux93_inw5),
.DataIn_6(MEMOCMux93_inw6),
.DataIn_7(MEMOCMux93_inw7),
.DataIn_8(MEMOCMux93_inw8),
.DataIn_9(MEMOCMux93_inw9),
.DataIn_10(MEMOCMux93_inw10),
.DataOut_1(MEMOCMux93_outw1),
.sel(MEMOCMux93_selw));
defparam MEMOCMux93.Mux_BW = 32;
assign MEMC93_data_from_Core = MEMOCMux93_outw1;
assign MEMOCMux93_inw1 = dataOutW[31:0]; 
assign MEMOCMux93_inw2 = dataOutW[63:32]; 
assign MEMOCMux93_inw3 = dataOutW[95:64]; 
assign MEMOCMux93_inw4 = dataOutW[127:96]; 
assign MEMOCMux93_inw5 = dataOutW[159:128]; 
assign MEMOCMux93_inw6 = dataOutW[191:160]; 
assign MEMOCMux93_inw7 = dataOutW[223:192]; 
assign MEMOCMux93_inw8 = dataOutW[255:224]; 
assign MEMOCMux93_inw9 = dataOutW[287:256]; 
assign MEMOCMux93_inw10 = globalDataIn[3007:2976]; 
assign MEMOCMux93_selw = mOutConfigW[375:372]; 
assign MEMC93_data_out_ctx2 = mDataFromMem[3007:2976]; 
assign mDataToMem[3007:2976] = MEMC93_data_in_ctx1; 
assign globalDataOut[3007:2976] = MEMC93_data_to_Core; 
assign MEMC93_valid_ctx1 = valid1[93:93]; 
assign MEMC93_write_en_ctx1 = WEn1[93:93]; 
assign MEMC93_stride_ctx1 = stride1[93:93]; 
assign MEMC93_start_addr_ctx1 = startAddr1[563:558]; 
assign MEMC93_burst_count_ctx1 = count1[657:651]; 
assign mAddr1[563:558] = MEMC93_addr_out_ctx1; 
assign mEn1[93:93] = MEMC93_mem_en_ctx1; 
assign mWEn1[93:93] = MEMC93_write_mem_en_ctx1; 
assign MEMC93_valid_ctx2 = valid2[93:93]; 
assign MEMC93_write_en_ctx2 = WEn2[93:93]; 
assign MEMC93_stride_ctx2 = stride2[93:93]; 
assign MEMC93_start_addr_ctx2 = startAddr2[563:558]; 
assign mAddr2[563:558] = MEMC93_addr_out_ctx2; 
assign MEMC93_burst_count_ctx2 = count2[657:651]; 
assign mEn2[93:93] = MEMC93_mem_en_ctx2; 
assign mWEn2[93:93] = MEMC93_write_mem_en_ctx2; 
wire [31:0] MEMOCMux94_inw1;
wire [31:0] MEMOCMux94_inw2;
wire [31:0] MEMOCMux94_inw3;
wire [31:0] MEMOCMux94_inw4;
wire [31:0] MEMOCMux94_inw5;
wire [31:0] MEMOCMux94_inw6;
wire [31:0] MEMOCMux94_inw7;
wire [31:0] MEMOCMux94_inw8;
wire [31:0] MEMOCMux94_inw9;
wire [31:0] MEMOCMux94_inw10;
wire [31:0] MEMOCMux94_outw1;
wire [3:0] MEMOCMux94_selw;
HA_10IM MEMOCMux94 (
.DataIn_1(MEMOCMux94_inw1),
.DataIn_2(MEMOCMux94_inw2),
.DataIn_3(MEMOCMux94_inw3),
.DataIn_4(MEMOCMux94_inw4),
.DataIn_5(MEMOCMux94_inw5),
.DataIn_6(MEMOCMux94_inw6),
.DataIn_7(MEMOCMux94_inw7),
.DataIn_8(MEMOCMux94_inw8),
.DataIn_9(MEMOCMux94_inw9),
.DataIn_10(MEMOCMux94_inw10),
.DataOut_1(MEMOCMux94_outw1),
.sel(MEMOCMux94_selw));
defparam MEMOCMux94.Mux_BW = 32;
assign MEMC94_data_from_Core = MEMOCMux94_outw1;
assign MEMOCMux94_inw1 = dataOutW[31:0]; 
assign MEMOCMux94_inw2 = dataOutW[63:32]; 
assign MEMOCMux94_inw3 = dataOutW[95:64]; 
assign MEMOCMux94_inw4 = dataOutW[127:96]; 
assign MEMOCMux94_inw5 = dataOutW[159:128]; 
assign MEMOCMux94_inw6 = dataOutW[191:160]; 
assign MEMOCMux94_inw7 = dataOutW[223:192]; 
assign MEMOCMux94_inw8 = dataOutW[255:224]; 
assign MEMOCMux94_inw9 = dataOutW[287:256]; 
assign MEMOCMux94_inw10 = globalDataIn[3039:3008]; 
assign MEMOCMux94_selw = mOutConfigW[379:376]; 
assign MEMC94_data_out_ctx2 = mDataFromMem[3039:3008]; 
assign mDataToMem[3039:3008] = MEMC94_data_in_ctx1; 
assign globalDataOut[3039:3008] = MEMC94_data_to_Core; 
assign MEMC94_valid_ctx1 = valid1[94:94]; 
assign MEMC94_write_en_ctx1 = WEn1[94:94]; 
assign MEMC94_stride_ctx1 = stride1[94:94]; 
assign MEMC94_start_addr_ctx1 = startAddr1[569:564]; 
assign MEMC94_burst_count_ctx1 = count1[664:658]; 
assign mAddr1[569:564] = MEMC94_addr_out_ctx1; 
assign mEn1[94:94] = MEMC94_mem_en_ctx1; 
assign mWEn1[94:94] = MEMC94_write_mem_en_ctx1; 
assign MEMC94_valid_ctx2 = valid2[94:94]; 
assign MEMC94_write_en_ctx2 = WEn2[94:94]; 
assign MEMC94_stride_ctx2 = stride2[94:94]; 
assign MEMC94_start_addr_ctx2 = startAddr2[569:564]; 
assign mAddr2[569:564] = MEMC94_addr_out_ctx2; 
assign MEMC94_burst_count_ctx2 = count2[664:658]; 
assign mEn2[94:94] = MEMC94_mem_en_ctx2; 
assign mWEn2[94:94] = MEMC94_write_mem_en_ctx2; 
wire [31:0] MEMOCMux95_inw1;
wire [31:0] MEMOCMux95_inw2;
wire [31:0] MEMOCMux95_inw3;
wire [31:0] MEMOCMux95_inw4;
wire [31:0] MEMOCMux95_inw5;
wire [31:0] MEMOCMux95_inw6;
wire [31:0] MEMOCMux95_inw7;
wire [31:0] MEMOCMux95_inw8;
wire [31:0] MEMOCMux95_inw9;
wire [31:0] MEMOCMux95_inw10;
wire [31:0] MEMOCMux95_outw1;
wire [3:0] MEMOCMux95_selw;
HA_10IM MEMOCMux95 (
.DataIn_1(MEMOCMux95_inw1),
.DataIn_2(MEMOCMux95_inw2),
.DataIn_3(MEMOCMux95_inw3),
.DataIn_4(MEMOCMux95_inw4),
.DataIn_5(MEMOCMux95_inw5),
.DataIn_6(MEMOCMux95_inw6),
.DataIn_7(MEMOCMux95_inw7),
.DataIn_8(MEMOCMux95_inw8),
.DataIn_9(MEMOCMux95_inw9),
.DataIn_10(MEMOCMux95_inw10),
.DataOut_1(MEMOCMux95_outw1),
.sel(MEMOCMux95_selw));
defparam MEMOCMux95.Mux_BW = 32;
assign MEMC95_data_from_Core = MEMOCMux95_outw1;
assign MEMOCMux95_inw1 = dataOutW[31:0]; 
assign MEMOCMux95_inw2 = dataOutW[63:32]; 
assign MEMOCMux95_inw3 = dataOutW[95:64]; 
assign MEMOCMux95_inw4 = dataOutW[127:96]; 
assign MEMOCMux95_inw5 = dataOutW[159:128]; 
assign MEMOCMux95_inw6 = dataOutW[191:160]; 
assign MEMOCMux95_inw7 = dataOutW[223:192]; 
assign MEMOCMux95_inw8 = dataOutW[255:224]; 
assign MEMOCMux95_inw9 = dataOutW[287:256]; 
assign MEMOCMux95_inw10 = globalDataIn[3071:3040]; 
assign MEMOCMux95_selw = mOutConfigW[383:380]; 
assign MEMC95_data_out_ctx2 = mDataFromMem[3071:3040]; 
assign mDataToMem[3071:3040] = MEMC95_data_in_ctx1; 
assign globalDataOut[3071:3040] = MEMC95_data_to_Core; 
assign MEMC95_valid_ctx1 = valid1[95:95]; 
assign MEMC95_write_en_ctx1 = WEn1[95:95]; 
assign MEMC95_stride_ctx1 = stride1[95:95]; 
assign MEMC95_start_addr_ctx1 = startAddr1[575:570]; 
assign MEMC95_burst_count_ctx1 = count1[671:665]; 
assign mAddr1[575:570] = MEMC95_addr_out_ctx1; 
assign mEn1[95:95] = MEMC95_mem_en_ctx1; 
assign mWEn1[95:95] = MEMC95_write_mem_en_ctx1; 
assign MEMC95_valid_ctx2 = valid2[95:95]; 
assign MEMC95_write_en_ctx2 = WEn2[95:95]; 
assign MEMC95_stride_ctx2 = stride2[95:95]; 
assign MEMC95_start_addr_ctx2 = startAddr2[575:570]; 
assign mAddr2[575:570] = MEMC95_addr_out_ctx2; 
assign MEMC95_burst_count_ctx2 = count2[671:665]; 
assign mEn2[95:95] = MEMC95_mem_en_ctx2; 
assign mWEn2[95:95] = MEMC95_write_mem_en_ctx2; 
wire [31:0] MEMOCMux96_inw1;
wire [31:0] MEMOCMux96_inw2;
wire [31:0] MEMOCMux96_inw3;
wire [31:0] MEMOCMux96_inw4;
wire [31:0] MEMOCMux96_inw5;
wire [31:0] MEMOCMux96_inw6;
wire [31:0] MEMOCMux96_inw7;
wire [31:0] MEMOCMux96_inw8;
wire [31:0] MEMOCMux96_inw9;
wire [31:0] MEMOCMux96_inw10;
wire [31:0] MEMOCMux96_outw1;
wire [3:0] MEMOCMux96_selw;
HA_10IM MEMOCMux96 (
.DataIn_1(MEMOCMux96_inw1),
.DataIn_2(MEMOCMux96_inw2),
.DataIn_3(MEMOCMux96_inw3),
.DataIn_4(MEMOCMux96_inw4),
.DataIn_5(MEMOCMux96_inw5),
.DataIn_6(MEMOCMux96_inw6),
.DataIn_7(MEMOCMux96_inw7),
.DataIn_8(MEMOCMux96_inw8),
.DataIn_9(MEMOCMux96_inw9),
.DataIn_10(MEMOCMux96_inw10),
.DataOut_1(MEMOCMux96_outw1),
.sel(MEMOCMux96_selw));
defparam MEMOCMux96.Mux_BW = 32;
assign MEMC96_data_from_Core = MEMOCMux96_outw1;
assign MEMOCMux96_inw1 = dataOutW[31:0]; 
assign MEMOCMux96_inw2 = dataOutW[63:32]; 
assign MEMOCMux96_inw3 = dataOutW[95:64]; 
assign MEMOCMux96_inw4 = dataOutW[127:96]; 
assign MEMOCMux96_inw5 = dataOutW[159:128]; 
assign MEMOCMux96_inw6 = dataOutW[191:160]; 
assign MEMOCMux96_inw7 = dataOutW[223:192]; 
assign MEMOCMux96_inw8 = dataOutW[255:224]; 
assign MEMOCMux96_inw9 = dataOutW[287:256]; 
assign MEMOCMux96_inw10 = globalDataIn[3103:3072]; 
assign MEMOCMux96_selw = mOutConfigW[387:384]; 
assign MEMC96_data_out_ctx2 = mDataFromMem[3103:3072]; 
assign mDataToMem[3103:3072] = MEMC96_data_in_ctx1; 
assign globalDataOut[3103:3072] = MEMC96_data_to_Core; 
assign MEMC96_valid_ctx1 = valid1[96:96]; 
assign MEMC96_write_en_ctx1 = WEn1[96:96]; 
assign MEMC96_stride_ctx1 = stride1[96:96]; 
assign MEMC96_start_addr_ctx1 = startAddr1[581:576]; 
assign MEMC96_burst_count_ctx1 = count1[678:672]; 
assign mAddr1[581:576] = MEMC96_addr_out_ctx1; 
assign mEn1[96:96] = MEMC96_mem_en_ctx1; 
assign mWEn1[96:96] = MEMC96_write_mem_en_ctx1; 
assign MEMC96_valid_ctx2 = valid2[96:96]; 
assign MEMC96_write_en_ctx2 = WEn2[96:96]; 
assign MEMC96_stride_ctx2 = stride2[96:96]; 
assign MEMC96_start_addr_ctx2 = startAddr2[581:576]; 
assign mAddr2[581:576] = MEMC96_addr_out_ctx2; 
assign MEMC96_burst_count_ctx2 = count2[678:672]; 
assign mEn2[96:96] = MEMC96_mem_en_ctx2; 
assign mWEn2[96:96] = MEMC96_write_mem_en_ctx2; 
wire [31:0] MEMOCMux97_inw1;
wire [31:0] MEMOCMux97_inw2;
wire [31:0] MEMOCMux97_inw3;
wire [31:0] MEMOCMux97_inw4;
wire [31:0] MEMOCMux97_inw5;
wire [31:0] MEMOCMux97_inw6;
wire [31:0] MEMOCMux97_inw7;
wire [31:0] MEMOCMux97_inw8;
wire [31:0] MEMOCMux97_inw9;
wire [31:0] MEMOCMux97_inw10;
wire [31:0] MEMOCMux97_outw1;
wire [3:0] MEMOCMux97_selw;
HA_10IM MEMOCMux97 (
.DataIn_1(MEMOCMux97_inw1),
.DataIn_2(MEMOCMux97_inw2),
.DataIn_3(MEMOCMux97_inw3),
.DataIn_4(MEMOCMux97_inw4),
.DataIn_5(MEMOCMux97_inw5),
.DataIn_6(MEMOCMux97_inw6),
.DataIn_7(MEMOCMux97_inw7),
.DataIn_8(MEMOCMux97_inw8),
.DataIn_9(MEMOCMux97_inw9),
.DataIn_10(MEMOCMux97_inw10),
.DataOut_1(MEMOCMux97_outw1),
.sel(MEMOCMux97_selw));
defparam MEMOCMux97.Mux_BW = 32;
assign MEMC97_data_from_Core = MEMOCMux97_outw1;
assign MEMOCMux97_inw1 = dataOutW[31:0]; 
assign MEMOCMux97_inw2 = dataOutW[63:32]; 
assign MEMOCMux97_inw3 = dataOutW[95:64]; 
assign MEMOCMux97_inw4 = dataOutW[127:96]; 
assign MEMOCMux97_inw5 = dataOutW[159:128]; 
assign MEMOCMux97_inw6 = dataOutW[191:160]; 
assign MEMOCMux97_inw7 = dataOutW[223:192]; 
assign MEMOCMux97_inw8 = dataOutW[255:224]; 
assign MEMOCMux97_inw9 = dataOutW[287:256]; 
assign MEMOCMux97_inw10 = globalDataIn[3135:3104]; 
assign MEMOCMux97_selw = mOutConfigW[391:388]; 
assign MEMC97_data_out_ctx2 = mDataFromMem[3135:3104]; 
assign mDataToMem[3135:3104] = MEMC97_data_in_ctx1; 
assign globalDataOut[3135:3104] = MEMC97_data_to_Core; 
assign MEMC97_valid_ctx1 = valid1[97:97]; 
assign MEMC97_write_en_ctx1 = WEn1[97:97]; 
assign MEMC97_stride_ctx1 = stride1[97:97]; 
assign MEMC97_start_addr_ctx1 = startAddr1[587:582]; 
assign MEMC97_burst_count_ctx1 = count1[685:679]; 
assign mAddr1[587:582] = MEMC97_addr_out_ctx1; 
assign mEn1[97:97] = MEMC97_mem_en_ctx1; 
assign mWEn1[97:97] = MEMC97_write_mem_en_ctx1; 
assign MEMC97_valid_ctx2 = valid2[97:97]; 
assign MEMC97_write_en_ctx2 = WEn2[97:97]; 
assign MEMC97_stride_ctx2 = stride2[97:97]; 
assign MEMC97_start_addr_ctx2 = startAddr2[587:582]; 
assign mAddr2[587:582] = MEMC97_addr_out_ctx2; 
assign MEMC97_burst_count_ctx2 = count2[685:679]; 
assign mEn2[97:97] = MEMC97_mem_en_ctx2; 
assign mWEn2[97:97] = MEMC97_write_mem_en_ctx2; 
wire [31:0] MEMOCMux98_inw1;
wire [31:0] MEMOCMux98_inw2;
wire [31:0] MEMOCMux98_inw3;
wire [31:0] MEMOCMux98_inw4;
wire [31:0] MEMOCMux98_inw5;
wire [31:0] MEMOCMux98_inw6;
wire [31:0] MEMOCMux98_inw7;
wire [31:0] MEMOCMux98_inw8;
wire [31:0] MEMOCMux98_inw9;
wire [31:0] MEMOCMux98_inw10;
wire [31:0] MEMOCMux98_outw1;
wire [3:0] MEMOCMux98_selw;
HA_10IM MEMOCMux98 (
.DataIn_1(MEMOCMux98_inw1),
.DataIn_2(MEMOCMux98_inw2),
.DataIn_3(MEMOCMux98_inw3),
.DataIn_4(MEMOCMux98_inw4),
.DataIn_5(MEMOCMux98_inw5),
.DataIn_6(MEMOCMux98_inw6),
.DataIn_7(MEMOCMux98_inw7),
.DataIn_8(MEMOCMux98_inw8),
.DataIn_9(MEMOCMux98_inw9),
.DataIn_10(MEMOCMux98_inw10),
.DataOut_1(MEMOCMux98_outw1),
.sel(MEMOCMux98_selw));
defparam MEMOCMux98.Mux_BW = 32;
assign MEMC98_data_from_Core = MEMOCMux98_outw1;
assign MEMOCMux98_inw1 = dataOutW[31:0]; 
assign MEMOCMux98_inw2 = dataOutW[63:32]; 
assign MEMOCMux98_inw3 = dataOutW[95:64]; 
assign MEMOCMux98_inw4 = dataOutW[127:96]; 
assign MEMOCMux98_inw5 = dataOutW[159:128]; 
assign MEMOCMux98_inw6 = dataOutW[191:160]; 
assign MEMOCMux98_inw7 = dataOutW[223:192]; 
assign MEMOCMux98_inw8 = dataOutW[255:224]; 
assign MEMOCMux98_inw9 = dataOutW[287:256]; 
assign MEMOCMux98_inw10 = globalDataIn[3167:3136]; 
assign MEMOCMux98_selw = mOutConfigW[395:392]; 
assign MEMC98_data_out_ctx2 = mDataFromMem[3167:3136]; 
assign mDataToMem[3167:3136] = MEMC98_data_in_ctx1; 
assign globalDataOut[3167:3136] = MEMC98_data_to_Core; 
assign MEMC98_valid_ctx1 = valid1[98:98]; 
assign MEMC98_write_en_ctx1 = WEn1[98:98]; 
assign MEMC98_stride_ctx1 = stride1[98:98]; 
assign MEMC98_start_addr_ctx1 = startAddr1[593:588]; 
assign MEMC98_burst_count_ctx1 = count1[692:686]; 
assign mAddr1[593:588] = MEMC98_addr_out_ctx1; 
assign mEn1[98:98] = MEMC98_mem_en_ctx1; 
assign mWEn1[98:98] = MEMC98_write_mem_en_ctx1; 
assign MEMC98_valid_ctx2 = valid2[98:98]; 
assign MEMC98_write_en_ctx2 = WEn2[98:98]; 
assign MEMC98_stride_ctx2 = stride2[98:98]; 
assign MEMC98_start_addr_ctx2 = startAddr2[593:588]; 
assign mAddr2[593:588] = MEMC98_addr_out_ctx2; 
assign MEMC98_burst_count_ctx2 = count2[692:686]; 
assign mEn2[98:98] = MEMC98_mem_en_ctx2; 
assign mWEn2[98:98] = MEMC98_write_mem_en_ctx2; 
wire [31:0] MEMOCMux99_inw1;
wire [31:0] MEMOCMux99_inw2;
wire [31:0] MEMOCMux99_inw3;
wire [31:0] MEMOCMux99_inw4;
wire [31:0] MEMOCMux99_inw5;
wire [31:0] MEMOCMux99_inw6;
wire [31:0] MEMOCMux99_inw7;
wire [31:0] MEMOCMux99_inw8;
wire [31:0] MEMOCMux99_inw9;
wire [31:0] MEMOCMux99_inw10;
wire [31:0] MEMOCMux99_outw1;
wire [3:0] MEMOCMux99_selw;
HA_10IM MEMOCMux99 (
.DataIn_1(MEMOCMux99_inw1),
.DataIn_2(MEMOCMux99_inw2),
.DataIn_3(MEMOCMux99_inw3),
.DataIn_4(MEMOCMux99_inw4),
.DataIn_5(MEMOCMux99_inw5),
.DataIn_6(MEMOCMux99_inw6),
.DataIn_7(MEMOCMux99_inw7),
.DataIn_8(MEMOCMux99_inw8),
.DataIn_9(MEMOCMux99_inw9),
.DataIn_10(MEMOCMux99_inw10),
.DataOut_1(MEMOCMux99_outw1),
.sel(MEMOCMux99_selw));
defparam MEMOCMux99.Mux_BW = 32;
assign MEMC99_data_from_Core = MEMOCMux99_outw1;
assign MEMOCMux99_inw1 = dataOutW[31:0]; 
assign MEMOCMux99_inw2 = dataOutW[63:32]; 
assign MEMOCMux99_inw3 = dataOutW[95:64]; 
assign MEMOCMux99_inw4 = dataOutW[127:96]; 
assign MEMOCMux99_inw5 = dataOutW[159:128]; 
assign MEMOCMux99_inw6 = dataOutW[191:160]; 
assign MEMOCMux99_inw7 = dataOutW[223:192]; 
assign MEMOCMux99_inw8 = dataOutW[255:224]; 
assign MEMOCMux99_inw9 = dataOutW[287:256]; 
assign MEMOCMux99_inw10 = globalDataIn[3199:3168]; 
assign MEMOCMux99_selw = mOutConfigW[399:396]; 
assign MEMC99_data_out_ctx2 = mDataFromMem[3199:3168]; 
assign mDataToMem[3199:3168] = MEMC99_data_in_ctx1; 
assign globalDataOut[3199:3168] = MEMC99_data_to_Core; 
assign MEMC99_valid_ctx1 = valid1[99:99]; 
assign MEMC99_write_en_ctx1 = WEn1[99:99]; 
assign MEMC99_stride_ctx1 = stride1[99:99]; 
assign MEMC99_start_addr_ctx1 = startAddr1[599:594]; 
assign MEMC99_burst_count_ctx1 = count1[699:693]; 
assign mAddr1[599:594] = MEMC99_addr_out_ctx1; 
assign mEn1[99:99] = MEMC99_mem_en_ctx1; 
assign mWEn1[99:99] = MEMC99_write_mem_en_ctx1; 
assign MEMC99_valid_ctx2 = valid2[99:99]; 
assign MEMC99_write_en_ctx2 = WEn2[99:99]; 
assign MEMC99_stride_ctx2 = stride2[99:99]; 
assign MEMC99_start_addr_ctx2 = startAddr2[599:594]; 
assign mAddr2[599:594] = MEMC99_addr_out_ctx2; 
assign MEMC99_burst_count_ctx2 = count2[699:693]; 
assign mEn2[99:99] = MEMC99_mem_en_ctx2; 
assign mWEn2[99:99] = MEMC99_write_mem_en_ctx2; 
wire [31:0] MEMOCMux100_inw1;
wire [31:0] MEMOCMux100_inw2;
wire [31:0] MEMOCMux100_inw3;
wire [31:0] MEMOCMux100_inw4;
wire [31:0] MEMOCMux100_inw5;
wire [31:0] MEMOCMux100_inw6;
wire [31:0] MEMOCMux100_inw7;
wire [31:0] MEMOCMux100_inw8;
wire [31:0] MEMOCMux100_inw9;
wire [31:0] MEMOCMux100_inw10;
wire [31:0] MEMOCMux100_outw1;
wire [3:0] MEMOCMux100_selw;
HA_10IM MEMOCMux100 (
.DataIn_1(MEMOCMux100_inw1),
.DataIn_2(MEMOCMux100_inw2),
.DataIn_3(MEMOCMux100_inw3),
.DataIn_4(MEMOCMux100_inw4),
.DataIn_5(MEMOCMux100_inw5),
.DataIn_6(MEMOCMux100_inw6),
.DataIn_7(MEMOCMux100_inw7),
.DataIn_8(MEMOCMux100_inw8),
.DataIn_9(MEMOCMux100_inw9),
.DataIn_10(MEMOCMux100_inw10),
.DataOut_1(MEMOCMux100_outw1),
.sel(MEMOCMux100_selw));
defparam MEMOCMux100.Mux_BW = 32;
assign MEMC100_data_from_Core = MEMOCMux100_outw1;
assign MEMOCMux100_inw1 = dataOutW[31:0]; 
assign MEMOCMux100_inw2 = dataOutW[63:32]; 
assign MEMOCMux100_inw3 = dataOutW[95:64]; 
assign MEMOCMux100_inw4 = dataOutW[127:96]; 
assign MEMOCMux100_inw5 = dataOutW[159:128]; 
assign MEMOCMux100_inw6 = dataOutW[191:160]; 
assign MEMOCMux100_inw7 = dataOutW[223:192]; 
assign MEMOCMux100_inw8 = dataOutW[255:224]; 
assign MEMOCMux100_inw9 = dataOutW[287:256]; 
assign MEMOCMux100_inw10 = globalDataIn[3231:3200]; 
assign MEMOCMux100_selw = mOutConfigW[403:400]; 
assign MEMC100_data_out_ctx2 = mDataFromMem[3231:3200]; 
assign mDataToMem[3231:3200] = MEMC100_data_in_ctx1; 
assign globalDataOut[3231:3200] = MEMC100_data_to_Core; 
assign MEMC100_valid_ctx1 = valid1[100:100]; 
assign MEMC100_write_en_ctx1 = WEn1[100:100]; 
assign MEMC100_stride_ctx1 = stride1[100:100]; 
assign MEMC100_start_addr_ctx1 = startAddr1[605:600]; 
assign MEMC100_burst_count_ctx1 = count1[706:700]; 
assign mAddr1[605:600] = MEMC100_addr_out_ctx1; 
assign mEn1[100:100] = MEMC100_mem_en_ctx1; 
assign mWEn1[100:100] = MEMC100_write_mem_en_ctx1; 
assign MEMC100_valid_ctx2 = valid2[100:100]; 
assign MEMC100_write_en_ctx2 = WEn2[100:100]; 
assign MEMC100_stride_ctx2 = stride2[100:100]; 
assign MEMC100_start_addr_ctx2 = startAddr2[605:600]; 
assign mAddr2[605:600] = MEMC100_addr_out_ctx2; 
assign MEMC100_burst_count_ctx2 = count2[706:700]; 
assign mEn2[100:100] = MEMC100_mem_en_ctx2; 
assign mWEn2[100:100] = MEMC100_write_mem_en_ctx2; 
wire [31:0] MEMOCMux101_inw1;
wire [31:0] MEMOCMux101_inw2;
wire [31:0] MEMOCMux101_inw3;
wire [31:0] MEMOCMux101_inw4;
wire [31:0] MEMOCMux101_inw5;
wire [31:0] MEMOCMux101_inw6;
wire [31:0] MEMOCMux101_inw7;
wire [31:0] MEMOCMux101_inw8;
wire [31:0] MEMOCMux101_inw9;
wire [31:0] MEMOCMux101_inw10;
wire [31:0] MEMOCMux101_outw1;
wire [3:0] MEMOCMux101_selw;
HA_10IM MEMOCMux101 (
.DataIn_1(MEMOCMux101_inw1),
.DataIn_2(MEMOCMux101_inw2),
.DataIn_3(MEMOCMux101_inw3),
.DataIn_4(MEMOCMux101_inw4),
.DataIn_5(MEMOCMux101_inw5),
.DataIn_6(MEMOCMux101_inw6),
.DataIn_7(MEMOCMux101_inw7),
.DataIn_8(MEMOCMux101_inw8),
.DataIn_9(MEMOCMux101_inw9),
.DataIn_10(MEMOCMux101_inw10),
.DataOut_1(MEMOCMux101_outw1),
.sel(MEMOCMux101_selw));
defparam MEMOCMux101.Mux_BW = 32;
assign MEMC101_data_from_Core = MEMOCMux101_outw1;
assign MEMOCMux101_inw1 = dataOutW[31:0]; 
assign MEMOCMux101_inw2 = dataOutW[63:32]; 
assign MEMOCMux101_inw3 = dataOutW[95:64]; 
assign MEMOCMux101_inw4 = dataOutW[127:96]; 
assign MEMOCMux101_inw5 = dataOutW[159:128]; 
assign MEMOCMux101_inw6 = dataOutW[191:160]; 
assign MEMOCMux101_inw7 = dataOutW[223:192]; 
assign MEMOCMux101_inw8 = dataOutW[255:224]; 
assign MEMOCMux101_inw9 = dataOutW[287:256]; 
assign MEMOCMux101_inw10 = globalDataIn[3263:3232]; 
assign MEMOCMux101_selw = mOutConfigW[407:404]; 
assign MEMC101_data_out_ctx2 = mDataFromMem[3263:3232]; 
assign mDataToMem[3263:3232] = MEMC101_data_in_ctx1; 
assign globalDataOut[3263:3232] = MEMC101_data_to_Core; 
assign MEMC101_valid_ctx1 = valid1[101:101]; 
assign MEMC101_write_en_ctx1 = WEn1[101:101]; 
assign MEMC101_stride_ctx1 = stride1[101:101]; 
assign MEMC101_start_addr_ctx1 = startAddr1[611:606]; 
assign MEMC101_burst_count_ctx1 = count1[713:707]; 
assign mAddr1[611:606] = MEMC101_addr_out_ctx1; 
assign mEn1[101:101] = MEMC101_mem_en_ctx1; 
assign mWEn1[101:101] = MEMC101_write_mem_en_ctx1; 
assign MEMC101_valid_ctx2 = valid2[101:101]; 
assign MEMC101_write_en_ctx2 = WEn2[101:101]; 
assign MEMC101_stride_ctx2 = stride2[101:101]; 
assign MEMC101_start_addr_ctx2 = startAddr2[611:606]; 
assign mAddr2[611:606] = MEMC101_addr_out_ctx2; 
assign MEMC101_burst_count_ctx2 = count2[713:707]; 
assign mEn2[101:101] = MEMC101_mem_en_ctx2; 
assign mWEn2[101:101] = MEMC101_write_mem_en_ctx2; 
wire [31:0] MEMOCMux102_inw1;
wire [31:0] MEMOCMux102_inw2;
wire [31:0] MEMOCMux102_inw3;
wire [31:0] MEMOCMux102_inw4;
wire [31:0] MEMOCMux102_inw5;
wire [31:0] MEMOCMux102_inw6;
wire [31:0] MEMOCMux102_inw7;
wire [31:0] MEMOCMux102_inw8;
wire [31:0] MEMOCMux102_inw9;
wire [31:0] MEMOCMux102_inw10;
wire [31:0] MEMOCMux102_outw1;
wire [3:0] MEMOCMux102_selw;
HA_10IM MEMOCMux102 (
.DataIn_1(MEMOCMux102_inw1),
.DataIn_2(MEMOCMux102_inw2),
.DataIn_3(MEMOCMux102_inw3),
.DataIn_4(MEMOCMux102_inw4),
.DataIn_5(MEMOCMux102_inw5),
.DataIn_6(MEMOCMux102_inw6),
.DataIn_7(MEMOCMux102_inw7),
.DataIn_8(MEMOCMux102_inw8),
.DataIn_9(MEMOCMux102_inw9),
.DataIn_10(MEMOCMux102_inw10),
.DataOut_1(MEMOCMux102_outw1),
.sel(MEMOCMux102_selw));
defparam MEMOCMux102.Mux_BW = 32;
assign MEMC102_data_from_Core = MEMOCMux102_outw1;
assign MEMOCMux102_inw1 = dataOutW[31:0]; 
assign MEMOCMux102_inw2 = dataOutW[63:32]; 
assign MEMOCMux102_inw3 = dataOutW[95:64]; 
assign MEMOCMux102_inw4 = dataOutW[127:96]; 
assign MEMOCMux102_inw5 = dataOutW[159:128]; 
assign MEMOCMux102_inw6 = dataOutW[191:160]; 
assign MEMOCMux102_inw7 = dataOutW[223:192]; 
assign MEMOCMux102_inw8 = dataOutW[255:224]; 
assign MEMOCMux102_inw9 = dataOutW[287:256]; 
assign MEMOCMux102_inw10 = globalDataIn[3295:3264]; 
assign MEMOCMux102_selw = mOutConfigW[411:408]; 
assign MEMC102_data_out_ctx2 = mDataFromMem[3295:3264]; 
assign mDataToMem[3295:3264] = MEMC102_data_in_ctx1; 
assign globalDataOut[3295:3264] = MEMC102_data_to_Core; 
assign MEMC102_valid_ctx1 = valid1[102:102]; 
assign MEMC102_write_en_ctx1 = WEn1[102:102]; 
assign MEMC102_stride_ctx1 = stride1[102:102]; 
assign MEMC102_start_addr_ctx1 = startAddr1[617:612]; 
assign MEMC102_burst_count_ctx1 = count1[720:714]; 
assign mAddr1[617:612] = MEMC102_addr_out_ctx1; 
assign mEn1[102:102] = MEMC102_mem_en_ctx1; 
assign mWEn1[102:102] = MEMC102_write_mem_en_ctx1; 
assign MEMC102_valid_ctx2 = valid2[102:102]; 
assign MEMC102_write_en_ctx2 = WEn2[102:102]; 
assign MEMC102_stride_ctx2 = stride2[102:102]; 
assign MEMC102_start_addr_ctx2 = startAddr2[617:612]; 
assign mAddr2[617:612] = MEMC102_addr_out_ctx2; 
assign MEMC102_burst_count_ctx2 = count2[720:714]; 
assign mEn2[102:102] = MEMC102_mem_en_ctx2; 
assign mWEn2[102:102] = MEMC102_write_mem_en_ctx2; 
wire [31:0] MEMOCMux103_inw1;
wire [31:0] MEMOCMux103_inw2;
wire [31:0] MEMOCMux103_inw3;
wire [31:0] MEMOCMux103_inw4;
wire [31:0] MEMOCMux103_inw5;
wire [31:0] MEMOCMux103_inw6;
wire [31:0] MEMOCMux103_inw7;
wire [31:0] MEMOCMux103_inw8;
wire [31:0] MEMOCMux103_inw9;
wire [31:0] MEMOCMux103_inw10;
wire [31:0] MEMOCMux103_outw1;
wire [3:0] MEMOCMux103_selw;
HA_10IM MEMOCMux103 (
.DataIn_1(MEMOCMux103_inw1),
.DataIn_2(MEMOCMux103_inw2),
.DataIn_3(MEMOCMux103_inw3),
.DataIn_4(MEMOCMux103_inw4),
.DataIn_5(MEMOCMux103_inw5),
.DataIn_6(MEMOCMux103_inw6),
.DataIn_7(MEMOCMux103_inw7),
.DataIn_8(MEMOCMux103_inw8),
.DataIn_9(MEMOCMux103_inw9),
.DataIn_10(MEMOCMux103_inw10),
.DataOut_1(MEMOCMux103_outw1),
.sel(MEMOCMux103_selw));
defparam MEMOCMux103.Mux_BW = 32;
assign MEMC103_data_from_Core = MEMOCMux103_outw1;
assign MEMOCMux103_inw1 = dataOutW[31:0]; 
assign MEMOCMux103_inw2 = dataOutW[63:32]; 
assign MEMOCMux103_inw3 = dataOutW[95:64]; 
assign MEMOCMux103_inw4 = dataOutW[127:96]; 
assign MEMOCMux103_inw5 = dataOutW[159:128]; 
assign MEMOCMux103_inw6 = dataOutW[191:160]; 
assign MEMOCMux103_inw7 = dataOutW[223:192]; 
assign MEMOCMux103_inw8 = dataOutW[255:224]; 
assign MEMOCMux103_inw9 = dataOutW[287:256]; 
assign MEMOCMux103_inw10 = globalDataIn[3327:3296]; 
assign MEMOCMux103_selw = mOutConfigW[415:412]; 
assign MEMC103_data_out_ctx2 = mDataFromMem[3327:3296]; 
assign mDataToMem[3327:3296] = MEMC103_data_in_ctx1; 
assign globalDataOut[3327:3296] = MEMC103_data_to_Core; 
assign MEMC103_valid_ctx1 = valid1[103:103]; 
assign MEMC103_write_en_ctx1 = WEn1[103:103]; 
assign MEMC103_stride_ctx1 = stride1[103:103]; 
assign MEMC103_start_addr_ctx1 = startAddr1[623:618]; 
assign MEMC103_burst_count_ctx1 = count1[727:721]; 
assign mAddr1[623:618] = MEMC103_addr_out_ctx1; 
assign mEn1[103:103] = MEMC103_mem_en_ctx1; 
assign mWEn1[103:103] = MEMC103_write_mem_en_ctx1; 
assign MEMC103_valid_ctx2 = valid2[103:103]; 
assign MEMC103_write_en_ctx2 = WEn2[103:103]; 
assign MEMC103_stride_ctx2 = stride2[103:103]; 
assign MEMC103_start_addr_ctx2 = startAddr2[623:618]; 
assign mAddr2[623:618] = MEMC103_addr_out_ctx2; 
assign MEMC103_burst_count_ctx2 = count2[727:721]; 
assign mEn2[103:103] = MEMC103_mem_en_ctx2; 
assign mWEn2[103:103] = MEMC103_write_mem_en_ctx2; 
wire [31:0] MEMOCMux104_inw1;
wire [31:0] MEMOCMux104_inw2;
wire [31:0] MEMOCMux104_inw3;
wire [31:0] MEMOCMux104_inw4;
wire [31:0] MEMOCMux104_inw5;
wire [31:0] MEMOCMux104_inw6;
wire [31:0] MEMOCMux104_inw7;
wire [31:0] MEMOCMux104_inw8;
wire [31:0] MEMOCMux104_inw9;
wire [31:0] MEMOCMux104_inw10;
wire [31:0] MEMOCMux104_outw1;
wire [3:0] MEMOCMux104_selw;
HA_10IM MEMOCMux104 (
.DataIn_1(MEMOCMux104_inw1),
.DataIn_2(MEMOCMux104_inw2),
.DataIn_3(MEMOCMux104_inw3),
.DataIn_4(MEMOCMux104_inw4),
.DataIn_5(MEMOCMux104_inw5),
.DataIn_6(MEMOCMux104_inw6),
.DataIn_7(MEMOCMux104_inw7),
.DataIn_8(MEMOCMux104_inw8),
.DataIn_9(MEMOCMux104_inw9),
.DataIn_10(MEMOCMux104_inw10),
.DataOut_1(MEMOCMux104_outw1),
.sel(MEMOCMux104_selw));
defparam MEMOCMux104.Mux_BW = 32;
assign MEMC104_data_from_Core = MEMOCMux104_outw1;
assign MEMOCMux104_inw1 = dataOutW[31:0]; 
assign MEMOCMux104_inw2 = dataOutW[63:32]; 
assign MEMOCMux104_inw3 = dataOutW[95:64]; 
assign MEMOCMux104_inw4 = dataOutW[127:96]; 
assign MEMOCMux104_inw5 = dataOutW[159:128]; 
assign MEMOCMux104_inw6 = dataOutW[191:160]; 
assign MEMOCMux104_inw7 = dataOutW[223:192]; 
assign MEMOCMux104_inw8 = dataOutW[255:224]; 
assign MEMOCMux104_inw9 = dataOutW[287:256]; 
assign MEMOCMux104_inw10 = globalDataIn[3359:3328]; 
assign MEMOCMux104_selw = mOutConfigW[419:416]; 
assign MEMC104_data_out_ctx2 = mDataFromMem[3359:3328]; 
assign mDataToMem[3359:3328] = MEMC104_data_in_ctx1; 
assign globalDataOut[3359:3328] = MEMC104_data_to_Core; 
assign MEMC104_valid_ctx1 = valid1[104:104]; 
assign MEMC104_write_en_ctx1 = WEn1[104:104]; 
assign MEMC104_stride_ctx1 = stride1[104:104]; 
assign MEMC104_start_addr_ctx1 = startAddr1[629:624]; 
assign MEMC104_burst_count_ctx1 = count1[734:728]; 
assign mAddr1[629:624] = MEMC104_addr_out_ctx1; 
assign mEn1[104:104] = MEMC104_mem_en_ctx1; 
assign mWEn1[104:104] = MEMC104_write_mem_en_ctx1; 
assign MEMC104_valid_ctx2 = valid2[104:104]; 
assign MEMC104_write_en_ctx2 = WEn2[104:104]; 
assign MEMC104_stride_ctx2 = stride2[104:104]; 
assign MEMC104_start_addr_ctx2 = startAddr2[629:624]; 
assign mAddr2[629:624] = MEMC104_addr_out_ctx2; 
assign MEMC104_burst_count_ctx2 = count2[734:728]; 
assign mEn2[104:104] = MEMC104_mem_en_ctx2; 
assign mWEn2[104:104] = MEMC104_write_mem_en_ctx2; 
wire [31:0] MEMOCMux105_inw1;
wire [31:0] MEMOCMux105_inw2;
wire [31:0] MEMOCMux105_inw3;
wire [31:0] MEMOCMux105_inw4;
wire [31:0] MEMOCMux105_inw5;
wire [31:0] MEMOCMux105_inw6;
wire [31:0] MEMOCMux105_inw7;
wire [31:0] MEMOCMux105_inw8;
wire [31:0] MEMOCMux105_inw9;
wire [31:0] MEMOCMux105_inw10;
wire [31:0] MEMOCMux105_outw1;
wire [3:0] MEMOCMux105_selw;
HA_10IM MEMOCMux105 (
.DataIn_1(MEMOCMux105_inw1),
.DataIn_2(MEMOCMux105_inw2),
.DataIn_3(MEMOCMux105_inw3),
.DataIn_4(MEMOCMux105_inw4),
.DataIn_5(MEMOCMux105_inw5),
.DataIn_6(MEMOCMux105_inw6),
.DataIn_7(MEMOCMux105_inw7),
.DataIn_8(MEMOCMux105_inw8),
.DataIn_9(MEMOCMux105_inw9),
.DataIn_10(MEMOCMux105_inw10),
.DataOut_1(MEMOCMux105_outw1),
.sel(MEMOCMux105_selw));
defparam MEMOCMux105.Mux_BW = 32;
assign MEMC105_data_from_Core = MEMOCMux105_outw1;
assign MEMOCMux105_inw1 = dataOutW[31:0]; 
assign MEMOCMux105_inw2 = dataOutW[63:32]; 
assign MEMOCMux105_inw3 = dataOutW[95:64]; 
assign MEMOCMux105_inw4 = dataOutW[127:96]; 
assign MEMOCMux105_inw5 = dataOutW[159:128]; 
assign MEMOCMux105_inw6 = dataOutW[191:160]; 
assign MEMOCMux105_inw7 = dataOutW[223:192]; 
assign MEMOCMux105_inw8 = dataOutW[255:224]; 
assign MEMOCMux105_inw9 = dataOutW[287:256]; 
assign MEMOCMux105_inw10 = globalDataIn[3391:3360]; 
assign MEMOCMux105_selw = mOutConfigW[423:420]; 
assign MEMC105_data_out_ctx2 = mDataFromMem[3391:3360]; 
assign mDataToMem[3391:3360] = MEMC105_data_in_ctx1; 
assign globalDataOut[3391:3360] = MEMC105_data_to_Core; 
assign MEMC105_valid_ctx1 = valid1[105:105]; 
assign MEMC105_write_en_ctx1 = WEn1[105:105]; 
assign MEMC105_stride_ctx1 = stride1[105:105]; 
assign MEMC105_start_addr_ctx1 = startAddr1[635:630]; 
assign MEMC105_burst_count_ctx1 = count1[741:735]; 
assign mAddr1[635:630] = MEMC105_addr_out_ctx1; 
assign mEn1[105:105] = MEMC105_mem_en_ctx1; 
assign mWEn1[105:105] = MEMC105_write_mem_en_ctx1; 
assign MEMC105_valid_ctx2 = valid2[105:105]; 
assign MEMC105_write_en_ctx2 = WEn2[105:105]; 
assign MEMC105_stride_ctx2 = stride2[105:105]; 
assign MEMC105_start_addr_ctx2 = startAddr2[635:630]; 
assign mAddr2[635:630] = MEMC105_addr_out_ctx2; 
assign MEMC105_burst_count_ctx2 = count2[741:735]; 
assign mEn2[105:105] = MEMC105_mem_en_ctx2; 
assign mWEn2[105:105] = MEMC105_write_mem_en_ctx2; 
wire [31:0] MEMOCMux106_inw1;
wire [31:0] MEMOCMux106_inw2;
wire [31:0] MEMOCMux106_inw3;
wire [31:0] MEMOCMux106_inw4;
wire [31:0] MEMOCMux106_inw5;
wire [31:0] MEMOCMux106_inw6;
wire [31:0] MEMOCMux106_inw7;
wire [31:0] MEMOCMux106_inw8;
wire [31:0] MEMOCMux106_inw9;
wire [31:0] MEMOCMux106_inw10;
wire [31:0] MEMOCMux106_outw1;
wire [3:0] MEMOCMux106_selw;
HA_10IM MEMOCMux106 (
.DataIn_1(MEMOCMux106_inw1),
.DataIn_2(MEMOCMux106_inw2),
.DataIn_3(MEMOCMux106_inw3),
.DataIn_4(MEMOCMux106_inw4),
.DataIn_5(MEMOCMux106_inw5),
.DataIn_6(MEMOCMux106_inw6),
.DataIn_7(MEMOCMux106_inw7),
.DataIn_8(MEMOCMux106_inw8),
.DataIn_9(MEMOCMux106_inw9),
.DataIn_10(MEMOCMux106_inw10),
.DataOut_1(MEMOCMux106_outw1),
.sel(MEMOCMux106_selw));
defparam MEMOCMux106.Mux_BW = 32;
assign MEMC106_data_from_Core = MEMOCMux106_outw1;
assign MEMOCMux106_inw1 = dataOutW[31:0]; 
assign MEMOCMux106_inw2 = dataOutW[63:32]; 
assign MEMOCMux106_inw3 = dataOutW[95:64]; 
assign MEMOCMux106_inw4 = dataOutW[127:96]; 
assign MEMOCMux106_inw5 = dataOutW[159:128]; 
assign MEMOCMux106_inw6 = dataOutW[191:160]; 
assign MEMOCMux106_inw7 = dataOutW[223:192]; 
assign MEMOCMux106_inw8 = dataOutW[255:224]; 
assign MEMOCMux106_inw9 = dataOutW[287:256]; 
assign MEMOCMux106_inw10 = globalDataIn[3423:3392]; 
assign MEMOCMux106_selw = mOutConfigW[427:424]; 
assign MEMC106_data_out_ctx2 = mDataFromMem[3423:3392]; 
assign mDataToMem[3423:3392] = MEMC106_data_in_ctx1; 
assign globalDataOut[3423:3392] = MEMC106_data_to_Core; 
assign MEMC106_valid_ctx1 = valid1[106:106]; 
assign MEMC106_write_en_ctx1 = WEn1[106:106]; 
assign MEMC106_stride_ctx1 = stride1[106:106]; 
assign MEMC106_start_addr_ctx1 = startAddr1[641:636]; 
assign MEMC106_burst_count_ctx1 = count1[748:742]; 
assign mAddr1[641:636] = MEMC106_addr_out_ctx1; 
assign mEn1[106:106] = MEMC106_mem_en_ctx1; 
assign mWEn1[106:106] = MEMC106_write_mem_en_ctx1; 
assign MEMC106_valid_ctx2 = valid2[106:106]; 
assign MEMC106_write_en_ctx2 = WEn2[106:106]; 
assign MEMC106_stride_ctx2 = stride2[106:106]; 
assign MEMC106_start_addr_ctx2 = startAddr2[641:636]; 
assign mAddr2[641:636] = MEMC106_addr_out_ctx2; 
assign MEMC106_burst_count_ctx2 = count2[748:742]; 
assign mEn2[106:106] = MEMC106_mem_en_ctx2; 
assign mWEn2[106:106] = MEMC106_write_mem_en_ctx2; 
wire [31:0] MEMOCMux107_inw1;
wire [31:0] MEMOCMux107_inw2;
wire [31:0] MEMOCMux107_inw3;
wire [31:0] MEMOCMux107_inw4;
wire [31:0] MEMOCMux107_inw5;
wire [31:0] MEMOCMux107_inw6;
wire [31:0] MEMOCMux107_inw7;
wire [31:0] MEMOCMux107_inw8;
wire [31:0] MEMOCMux107_inw9;
wire [31:0] MEMOCMux107_inw10;
wire [31:0] MEMOCMux107_outw1;
wire [3:0] MEMOCMux107_selw;
HA_10IM MEMOCMux107 (
.DataIn_1(MEMOCMux107_inw1),
.DataIn_2(MEMOCMux107_inw2),
.DataIn_3(MEMOCMux107_inw3),
.DataIn_4(MEMOCMux107_inw4),
.DataIn_5(MEMOCMux107_inw5),
.DataIn_6(MEMOCMux107_inw6),
.DataIn_7(MEMOCMux107_inw7),
.DataIn_8(MEMOCMux107_inw8),
.DataIn_9(MEMOCMux107_inw9),
.DataIn_10(MEMOCMux107_inw10),
.DataOut_1(MEMOCMux107_outw1),
.sel(MEMOCMux107_selw));
defparam MEMOCMux107.Mux_BW = 32;
assign MEMC107_data_from_Core = MEMOCMux107_outw1;
assign MEMOCMux107_inw1 = dataOutW[31:0]; 
assign MEMOCMux107_inw2 = dataOutW[63:32]; 
assign MEMOCMux107_inw3 = dataOutW[95:64]; 
assign MEMOCMux107_inw4 = dataOutW[127:96]; 
assign MEMOCMux107_inw5 = dataOutW[159:128]; 
assign MEMOCMux107_inw6 = dataOutW[191:160]; 
assign MEMOCMux107_inw7 = dataOutW[223:192]; 
assign MEMOCMux107_inw8 = dataOutW[255:224]; 
assign MEMOCMux107_inw9 = dataOutW[287:256]; 
assign MEMOCMux107_inw10 = globalDataIn[3455:3424]; 
assign MEMOCMux107_selw = mOutConfigW[431:428]; 
assign MEMC107_data_out_ctx2 = mDataFromMem[3455:3424]; 
assign mDataToMem[3455:3424] = MEMC107_data_in_ctx1; 
assign globalDataOut[3455:3424] = MEMC107_data_to_Core; 
assign MEMC107_valid_ctx1 = valid1[107:107]; 
assign MEMC107_write_en_ctx1 = WEn1[107:107]; 
assign MEMC107_stride_ctx1 = stride1[107:107]; 
assign MEMC107_start_addr_ctx1 = startAddr1[647:642]; 
assign MEMC107_burst_count_ctx1 = count1[755:749]; 
assign mAddr1[647:642] = MEMC107_addr_out_ctx1; 
assign mEn1[107:107] = MEMC107_mem_en_ctx1; 
assign mWEn1[107:107] = MEMC107_write_mem_en_ctx1; 
assign MEMC107_valid_ctx2 = valid2[107:107]; 
assign MEMC107_write_en_ctx2 = WEn2[107:107]; 
assign MEMC107_stride_ctx2 = stride2[107:107]; 
assign MEMC107_start_addr_ctx2 = startAddr2[647:642]; 
assign mAddr2[647:642] = MEMC107_addr_out_ctx2; 
assign MEMC107_burst_count_ctx2 = count2[755:749]; 
assign mEn2[107:107] = MEMC107_mem_en_ctx2; 
assign mWEn2[107:107] = MEMC107_write_mem_en_ctx2; 
assign dataInW[31:0] = MEMC0_data_to_Core; 
assign dataInW[63:32] = MEMC1_data_to_Core; 
assign dataInW[95:64] = MEMC2_data_to_Core; 
assign dataInW[127:96] = MEMC3_data_to_Core; 
assign dataInW[159:128] = MEMC4_data_to_Core; 
assign dataInW[191:160] = MEMC5_data_to_Core; 
assign dataInW[223:192] = MEMC6_data_to_Core; 
assign dataInW[255:224] = MEMC7_data_to_Core; 
assign dataInW[287:256] = MEMC8_data_to_Core; 
assign dataInW[319:288] = MEMC9_data_to_Core; 
assign dataInW[351:320] = MEMC10_data_to_Core; 
assign dataInW[383:352] = MEMC11_data_to_Core; 
assign dataInW[415:384] = MEMC12_data_to_Core; 
assign dataInW[447:416] = MEMC13_data_to_Core; 
assign dataInW[479:448] = MEMC14_data_to_Core; 
assign dataInW[511:480] = MEMC15_data_to_Core; 
assign dataInW[543:512] = MEMC16_data_to_Core; 
assign dataInW[575:544] = MEMC17_data_to_Core; 
assign dataInW[607:576] = MEMC18_data_to_Core; 
assign dataInW[639:608] = MEMC19_data_to_Core; 
assign dataInW[671:640] = MEMC20_data_to_Core; 
assign dataInW[703:672] = MEMC21_data_to_Core; 
assign dataInW[735:704] = MEMC22_data_to_Core; 
assign dataInW[767:736] = MEMC23_data_to_Core; 
assign dataInW[799:768] = MEMC24_data_to_Core; 
assign dataInW[831:800] = MEMC25_data_to_Core; 
assign dataInW[863:832] = MEMC26_data_to_Core; 
assign dataInW[895:864] = MEMC27_data_to_Core; 
assign dataInW[927:896] = MEMC28_data_to_Core; 
assign dataInW[959:928] = MEMC29_data_to_Core; 
assign dataInW[991:960] = MEMC30_data_to_Core; 
assign dataInW[1023:992] = MEMC31_data_to_Core; 
assign dataInW[1055:1024] = MEMC32_data_to_Core; 
assign dataInW[1087:1056] = MEMC33_data_to_Core; 
assign dataInW[1119:1088] = MEMC34_data_to_Core; 
assign dataInW[1151:1120] = MEMC35_data_to_Core; 
assign dataInW[1183:1152] = MEMC36_data_to_Core; 
assign dataInW[1215:1184] = MEMC37_data_to_Core; 
assign dataInW[1247:1216] = MEMC38_data_to_Core; 
assign dataInW[1279:1248] = MEMC39_data_to_Core; 
assign dataInW[1311:1280] = MEMC40_data_to_Core; 
assign dataInW[1343:1312] = MEMC41_data_to_Core; 
assign dataInW[1375:1344] = MEMC42_data_to_Core; 
assign dataInW[1407:1376] = MEMC43_data_to_Core; 
assign dataInW[1439:1408] = MEMC44_data_to_Core; 
assign dataInW[1471:1440] = MEMC45_data_to_Core; 
assign dataInW[1503:1472] = MEMC46_data_to_Core; 
assign dataInW[1535:1504] = MEMC47_data_to_Core; 
assign dataInW[1567:1536] = MEMC48_data_to_Core; 
assign dataInW[1599:1568] = MEMC49_data_to_Core; 
assign dataInW[1631:1600] = MEMC50_data_to_Core; 
assign dataInW[1663:1632] = MEMC51_data_to_Core; 
assign dataInW[1695:1664] = MEMC52_data_to_Core; 
assign dataInW[1727:1696] = MEMC53_data_to_Core; 
assign dataInW[1759:1728] = MEMC54_data_to_Core; 
assign dataInW[1791:1760] = MEMC55_data_to_Core; 
assign dataInW[1823:1792] = MEMC56_data_to_Core; 
assign dataInW[1855:1824] = MEMC57_data_to_Core; 
assign dataInW[1887:1856] = MEMC58_data_to_Core; 
assign dataInW[1919:1888] = MEMC59_data_to_Core; 
assign dataInW[1951:1920] = MEMC60_data_to_Core; 
assign dataInW[1983:1952] = MEMC61_data_to_Core; 
assign dataInW[2015:1984] = MEMC62_data_to_Core; 
assign dataInW[2047:2016] = MEMC63_data_to_Core; 
assign dataInW[2079:2048] = MEMC64_data_to_Core; 
assign dataInW[2111:2080] = MEMC65_data_to_Core; 
assign dataInW[2143:2112] = MEMC66_data_to_Core; 
assign dataInW[2175:2144] = MEMC67_data_to_Core; 
assign dataInW[2207:2176] = MEMC68_data_to_Core; 
assign dataInW[2239:2208] = MEMC69_data_to_Core; 
assign dataInW[2271:2240] = MEMC70_data_to_Core; 
assign dataInW[2303:2272] = MEMC71_data_to_Core; 
assign dataInW[2335:2304] = MEMC72_data_to_Core; 
assign dataInW[2367:2336] = MEMC73_data_to_Core; 
assign dataInW[2399:2368] = MEMC74_data_to_Core; 
assign dataInW[2431:2400] = MEMC75_data_to_Core; 
assign dataInW[2463:2432] = MEMC76_data_to_Core; 
assign dataInW[2495:2464] = MEMC77_data_to_Core; 
assign dataInW[2527:2496] = MEMC78_data_to_Core; 
assign dataInW[2559:2528] = MEMC79_data_to_Core; 
assign dataInW[2591:2560] = MEMC80_data_to_Core; 
assign dataInW[2623:2592] = MEMC81_data_to_Core; 
assign dataInW[2655:2624] = MEMC82_data_to_Core; 
assign dataInW[2687:2656] = MEMC83_data_to_Core; 
assign dataInW[2719:2688] = MEMC84_data_to_Core; 
assign dataInW[2751:2720] = MEMC85_data_to_Core; 
assign dataInW[2783:2752] = MEMC86_data_to_Core; 
assign dataInW[2815:2784] = MEMC87_data_to_Core; 
assign dataInW[2847:2816] = MEMC88_data_to_Core; 
assign dataInW[2879:2848] = MEMC89_data_to_Core; 
assign dataInW[2911:2880] = MEMC90_data_to_Core; 
assign dataInW[2943:2912] = MEMC91_data_to_Core; 
assign dataInW[2975:2944] = MEMC92_data_to_Core; 
assign dataInW[3007:2976] = MEMC93_data_to_Core; 
assign dataInW[3039:3008] = MEMC94_data_to_Core; 
assign dataInW[3071:3040] = MEMC95_data_to_Core; 
assign dataInW[3103:3072] = MEMC96_data_to_Core; 
assign dataInW[3135:3104] = MEMC97_data_to_Core; 
assign dataInW[3167:3136] = MEMC98_data_to_Core; 
assign dataInW[3199:3168] = MEMC99_data_to_Core; 
assign dataInW[3231:3200] = MEMC100_data_to_Core; 
assign dataInW[3263:3232] = MEMC101_data_to_Core; 
assign dataInW[3295:3264] = MEMC102_data_to_Core; 
assign dataInW[3327:3296] = MEMC103_data_to_Core; 
assign dataInW[3359:3328] = MEMC104_data_to_Core; 
assign dataInW[3391:3360] = MEMC105_data_to_Core; 
assign dataInW[3423:3392] = MEMC106_data_to_Core; 
assign dataInW[3455:3424] = MEMC107_data_to_Core; 
assign IMEMC_data_out_ctx2 = mIDataFromMem; 
assign mIDataToMem = IMEMC_data_in_ctx1; 
assign totalConfigInW = IMEMC_data_to_Core; 
assign IglobalDataOut = IMEMC_data_to_Core; 
assign IMEMC_data_from_Core = IglobalDataIn; 
assign IMEMC_valid_ctx1 = Ivalid1; 
assign IMEMC_write_en_ctx1 = IWEn1; 
assign IMEMC_stride_ctx1 = Istride1; 
assign IMEMC_start_addr_ctx1 = IstartAddr1; 
assign IMEMC_burst_count_ctx1 = Icount1; 
assign mIAddr1 = IMEMC_addr_out_ctx1; 
assign mIEn1 = IMEMC_mem_en_ctx1; 
assign mIWEn1 = IMEMC_write_mem_en_ctx1; 
assign IMEMC_valid_ctx2 = Ivalid2; 
assign IMEMC_write_en_ctx2 = IWEn2; 
assign IMEMC_stride_ctx2 = Istride2; 
assign IMEMC_start_addr_ctx2 = IstartAddr2; 
assign IMEMC_burst_count_ctx2 = Icount2; 
assign mIAddr2 = IMEMC_addr_out_ctx2; 
assign mIEn2 = IMEMC_mem_en_ctx2; 
assign mIWEn2 = IMEMC_write_mem_en_ctx2; 
endmodule
module MEMDock( mLocalDataIn, mLocalDataOut, mILocalDataIn, mILocalDataOut, MEMEnIn1, MEMRWEnIn1, MEMAddrIn1, IMEMEnIn1, IMEMRWEnIn1, IMEMAddrIn1, IMEMEnOut1, IMEMRWEnOut1, IMEMAddrOut1, MEMEnIn2, MEMRWEnIn2, MEMAddrIn2, IMEMEnIn2, IMEMRWEnIn2, IMEMAddrIn2, IMEMEnOut2, IMEMRWEnOut2, IMEMAddrOut2
,IMEMDataOut,IMEMDataIn
,MEMEnOut10,MEMDataOut0,MEMDataIn0,MEMAddrOut10,MEMRWEnOut10
,MEMEnOut20,MEMAddrOut20,MEMRWEnOut20
,MEMEnOut11,MEMDataOut1,MEMDataIn1,MEMAddrOut11,MEMRWEnOut11
,MEMEnOut21,MEMAddrOut21,MEMRWEnOut21
,MEMEnOut12,MEMDataOut2,MEMDataIn2,MEMAddrOut12,MEMRWEnOut12
,MEMEnOut22,MEMAddrOut22,MEMRWEnOut22
,MEMEnOut13,MEMDataOut3,MEMDataIn3,MEMAddrOut13,MEMRWEnOut13
,MEMEnOut23,MEMAddrOut23,MEMRWEnOut23
,MEMEnOut14,MEMDataOut4,MEMDataIn4,MEMAddrOut14,MEMRWEnOut14
,MEMEnOut24,MEMAddrOut24,MEMRWEnOut24
,MEMEnOut15,MEMDataOut5,MEMDataIn5,MEMAddrOut15,MEMRWEnOut15
,MEMEnOut25,MEMAddrOut25,MEMRWEnOut25
,MEMEnOut16,MEMDataOut6,MEMDataIn6,MEMAddrOut16,MEMRWEnOut16
,MEMEnOut26,MEMAddrOut26,MEMRWEnOut26
,MEMEnOut17,MEMDataOut7,MEMDataIn7,MEMAddrOut17,MEMRWEnOut17
,MEMEnOut27,MEMAddrOut27,MEMRWEnOut27
,MEMEnOut18,MEMDataOut8,MEMDataIn8,MEMAddrOut18,MEMRWEnOut18
,MEMEnOut28,MEMAddrOut28,MEMRWEnOut28
,MEMEnOut19,MEMDataOut9,MEMDataIn9,MEMAddrOut19,MEMRWEnOut19
,MEMEnOut29,MEMAddrOut29,MEMRWEnOut29
,MEMEnOut110,MEMDataOut10,MEMDataIn10,MEMAddrOut110,MEMRWEnOut110
,MEMEnOut210,MEMAddrOut210,MEMRWEnOut210
,MEMEnOut111,MEMDataOut11,MEMDataIn11,MEMAddrOut111,MEMRWEnOut111
,MEMEnOut211,MEMAddrOut211,MEMRWEnOut211
,MEMEnOut112,MEMDataOut12,MEMDataIn12,MEMAddrOut112,MEMRWEnOut112
,MEMEnOut212,MEMAddrOut212,MEMRWEnOut212
,MEMEnOut113,MEMDataOut13,MEMDataIn13,MEMAddrOut113,MEMRWEnOut113
,MEMEnOut213,MEMAddrOut213,MEMRWEnOut213
,MEMEnOut114,MEMDataOut14,MEMDataIn14,MEMAddrOut114,MEMRWEnOut114
,MEMEnOut214,MEMAddrOut214,MEMRWEnOut214
,MEMEnOut115,MEMDataOut15,MEMDataIn15,MEMAddrOut115,MEMRWEnOut115
,MEMEnOut215,MEMAddrOut215,MEMRWEnOut215
,MEMEnOut116,MEMDataOut16,MEMDataIn16,MEMAddrOut116,MEMRWEnOut116
,MEMEnOut216,MEMAddrOut216,MEMRWEnOut216
,MEMEnOut117,MEMDataOut17,MEMDataIn17,MEMAddrOut117,MEMRWEnOut117
,MEMEnOut217,MEMAddrOut217,MEMRWEnOut217
,MEMEnOut118,MEMDataOut18,MEMDataIn18,MEMAddrOut118,MEMRWEnOut118
,MEMEnOut218,MEMAddrOut218,MEMRWEnOut218
,MEMEnOut119,MEMDataOut19,MEMDataIn19,MEMAddrOut119,MEMRWEnOut119
,MEMEnOut219,MEMAddrOut219,MEMRWEnOut219
,MEMEnOut120,MEMDataOut20,MEMDataIn20,MEMAddrOut120,MEMRWEnOut120
,MEMEnOut220,MEMAddrOut220,MEMRWEnOut220
,MEMEnOut121,MEMDataOut21,MEMDataIn21,MEMAddrOut121,MEMRWEnOut121
,MEMEnOut221,MEMAddrOut221,MEMRWEnOut221
,MEMEnOut122,MEMDataOut22,MEMDataIn22,MEMAddrOut122,MEMRWEnOut122
,MEMEnOut222,MEMAddrOut222,MEMRWEnOut222
,MEMEnOut123,MEMDataOut23,MEMDataIn23,MEMAddrOut123,MEMRWEnOut123
,MEMEnOut223,MEMAddrOut223,MEMRWEnOut223
,MEMEnOut124,MEMDataOut24,MEMDataIn24,MEMAddrOut124,MEMRWEnOut124
,MEMEnOut224,MEMAddrOut224,MEMRWEnOut224
,MEMEnOut125,MEMDataOut25,MEMDataIn25,MEMAddrOut125,MEMRWEnOut125
,MEMEnOut225,MEMAddrOut225,MEMRWEnOut225
,MEMEnOut126,MEMDataOut26,MEMDataIn26,MEMAddrOut126,MEMRWEnOut126
,MEMEnOut226,MEMAddrOut226,MEMRWEnOut226
,MEMEnOut127,MEMDataOut27,MEMDataIn27,MEMAddrOut127,MEMRWEnOut127
,MEMEnOut227,MEMAddrOut227,MEMRWEnOut227
,MEMEnOut128,MEMDataOut28,MEMDataIn28,MEMAddrOut128,MEMRWEnOut128
,MEMEnOut228,MEMAddrOut228,MEMRWEnOut228
,MEMEnOut129,MEMDataOut29,MEMDataIn29,MEMAddrOut129,MEMRWEnOut129
,MEMEnOut229,MEMAddrOut229,MEMRWEnOut229
,MEMEnOut130,MEMDataOut30,MEMDataIn30,MEMAddrOut130,MEMRWEnOut130
,MEMEnOut230,MEMAddrOut230,MEMRWEnOut230
,MEMEnOut131,MEMDataOut31,MEMDataIn31,MEMAddrOut131,MEMRWEnOut131
,MEMEnOut231,MEMAddrOut231,MEMRWEnOut231
,MEMEnOut132,MEMDataOut32,MEMDataIn32,MEMAddrOut132,MEMRWEnOut132
,MEMEnOut232,MEMAddrOut232,MEMRWEnOut232
,MEMEnOut133,MEMDataOut33,MEMDataIn33,MEMAddrOut133,MEMRWEnOut133
,MEMEnOut233,MEMAddrOut233,MEMRWEnOut233
,MEMEnOut134,MEMDataOut34,MEMDataIn34,MEMAddrOut134,MEMRWEnOut134
,MEMEnOut234,MEMAddrOut234,MEMRWEnOut234
,MEMEnOut135,MEMDataOut35,MEMDataIn35,MEMAddrOut135,MEMRWEnOut135
,MEMEnOut235,MEMAddrOut235,MEMRWEnOut235
,MEMEnOut136,MEMDataOut36,MEMDataIn36,MEMAddrOut136,MEMRWEnOut136
,MEMEnOut236,MEMAddrOut236,MEMRWEnOut236
,MEMEnOut137,MEMDataOut37,MEMDataIn37,MEMAddrOut137,MEMRWEnOut137
,MEMEnOut237,MEMAddrOut237,MEMRWEnOut237
,MEMEnOut138,MEMDataOut38,MEMDataIn38,MEMAddrOut138,MEMRWEnOut138
,MEMEnOut238,MEMAddrOut238,MEMRWEnOut238
,MEMEnOut139,MEMDataOut39,MEMDataIn39,MEMAddrOut139,MEMRWEnOut139
,MEMEnOut239,MEMAddrOut239,MEMRWEnOut239
,MEMEnOut140,MEMDataOut40,MEMDataIn40,MEMAddrOut140,MEMRWEnOut140
,MEMEnOut240,MEMAddrOut240,MEMRWEnOut240
,MEMEnOut141,MEMDataOut41,MEMDataIn41,MEMAddrOut141,MEMRWEnOut141
,MEMEnOut241,MEMAddrOut241,MEMRWEnOut241
,MEMEnOut142,MEMDataOut42,MEMDataIn42,MEMAddrOut142,MEMRWEnOut142
,MEMEnOut242,MEMAddrOut242,MEMRWEnOut242
,MEMEnOut143,MEMDataOut43,MEMDataIn43,MEMAddrOut143,MEMRWEnOut143
,MEMEnOut243,MEMAddrOut243,MEMRWEnOut243
,MEMEnOut144,MEMDataOut44,MEMDataIn44,MEMAddrOut144,MEMRWEnOut144
,MEMEnOut244,MEMAddrOut244,MEMRWEnOut244
,MEMEnOut145,MEMDataOut45,MEMDataIn45,MEMAddrOut145,MEMRWEnOut145
,MEMEnOut245,MEMAddrOut245,MEMRWEnOut245
,MEMEnOut146,MEMDataOut46,MEMDataIn46,MEMAddrOut146,MEMRWEnOut146
,MEMEnOut246,MEMAddrOut246,MEMRWEnOut246
,MEMEnOut147,MEMDataOut47,MEMDataIn47,MEMAddrOut147,MEMRWEnOut147
,MEMEnOut247,MEMAddrOut247,MEMRWEnOut247
,MEMEnOut148,MEMDataOut48,MEMDataIn48,MEMAddrOut148,MEMRWEnOut148
,MEMEnOut248,MEMAddrOut248,MEMRWEnOut248
,MEMEnOut149,MEMDataOut49,MEMDataIn49,MEMAddrOut149,MEMRWEnOut149
,MEMEnOut249,MEMAddrOut249,MEMRWEnOut249
,MEMEnOut150,MEMDataOut50,MEMDataIn50,MEMAddrOut150,MEMRWEnOut150
,MEMEnOut250,MEMAddrOut250,MEMRWEnOut250
,MEMEnOut151,MEMDataOut51,MEMDataIn51,MEMAddrOut151,MEMRWEnOut151
,MEMEnOut251,MEMAddrOut251,MEMRWEnOut251
,MEMEnOut152,MEMDataOut52,MEMDataIn52,MEMAddrOut152,MEMRWEnOut152
,MEMEnOut252,MEMAddrOut252,MEMRWEnOut252
,MEMEnOut153,MEMDataOut53,MEMDataIn53,MEMAddrOut153,MEMRWEnOut153
,MEMEnOut253,MEMAddrOut253,MEMRWEnOut253
,MEMEnOut154,MEMDataOut54,MEMDataIn54,MEMAddrOut154,MEMRWEnOut154
,MEMEnOut254,MEMAddrOut254,MEMRWEnOut254
,MEMEnOut155,MEMDataOut55,MEMDataIn55,MEMAddrOut155,MEMRWEnOut155
,MEMEnOut255,MEMAddrOut255,MEMRWEnOut255
,MEMEnOut156,MEMDataOut56,MEMDataIn56,MEMAddrOut156,MEMRWEnOut156
,MEMEnOut256,MEMAddrOut256,MEMRWEnOut256
,MEMEnOut157,MEMDataOut57,MEMDataIn57,MEMAddrOut157,MEMRWEnOut157
,MEMEnOut257,MEMAddrOut257,MEMRWEnOut257
,MEMEnOut158,MEMDataOut58,MEMDataIn58,MEMAddrOut158,MEMRWEnOut158
,MEMEnOut258,MEMAddrOut258,MEMRWEnOut258
,MEMEnOut159,MEMDataOut59,MEMDataIn59,MEMAddrOut159,MEMRWEnOut159
,MEMEnOut259,MEMAddrOut259,MEMRWEnOut259
,MEMEnOut160,MEMDataOut60,MEMDataIn60,MEMAddrOut160,MEMRWEnOut160
,MEMEnOut260,MEMAddrOut260,MEMRWEnOut260
,MEMEnOut161,MEMDataOut61,MEMDataIn61,MEMAddrOut161,MEMRWEnOut161
,MEMEnOut261,MEMAddrOut261,MEMRWEnOut261
,MEMEnOut162,MEMDataOut62,MEMDataIn62,MEMAddrOut162,MEMRWEnOut162
,MEMEnOut262,MEMAddrOut262,MEMRWEnOut262
,MEMEnOut163,MEMDataOut63,MEMDataIn63,MEMAddrOut163,MEMRWEnOut163
,MEMEnOut263,MEMAddrOut263,MEMRWEnOut263
,MEMEnOut164,MEMDataOut64,MEMDataIn64,MEMAddrOut164,MEMRWEnOut164
,MEMEnOut264,MEMAddrOut264,MEMRWEnOut264
,MEMEnOut165,MEMDataOut65,MEMDataIn65,MEMAddrOut165,MEMRWEnOut165
,MEMEnOut265,MEMAddrOut265,MEMRWEnOut265
,MEMEnOut166,MEMDataOut66,MEMDataIn66,MEMAddrOut166,MEMRWEnOut166
,MEMEnOut266,MEMAddrOut266,MEMRWEnOut266
,MEMEnOut167,MEMDataOut67,MEMDataIn67,MEMAddrOut167,MEMRWEnOut167
,MEMEnOut267,MEMAddrOut267,MEMRWEnOut267
,MEMEnOut168,MEMDataOut68,MEMDataIn68,MEMAddrOut168,MEMRWEnOut168
,MEMEnOut268,MEMAddrOut268,MEMRWEnOut268
,MEMEnOut169,MEMDataOut69,MEMDataIn69,MEMAddrOut169,MEMRWEnOut169
,MEMEnOut269,MEMAddrOut269,MEMRWEnOut269
,MEMEnOut170,MEMDataOut70,MEMDataIn70,MEMAddrOut170,MEMRWEnOut170
,MEMEnOut270,MEMAddrOut270,MEMRWEnOut270
,MEMEnOut171,MEMDataOut71,MEMDataIn71,MEMAddrOut171,MEMRWEnOut171
,MEMEnOut271,MEMAddrOut271,MEMRWEnOut271
,MEMEnOut172,MEMDataOut72,MEMDataIn72,MEMAddrOut172,MEMRWEnOut172
,MEMEnOut272,MEMAddrOut272,MEMRWEnOut272
,MEMEnOut173,MEMDataOut73,MEMDataIn73,MEMAddrOut173,MEMRWEnOut173
,MEMEnOut273,MEMAddrOut273,MEMRWEnOut273
,MEMEnOut174,MEMDataOut74,MEMDataIn74,MEMAddrOut174,MEMRWEnOut174
,MEMEnOut274,MEMAddrOut274,MEMRWEnOut274
,MEMEnOut175,MEMDataOut75,MEMDataIn75,MEMAddrOut175,MEMRWEnOut175
,MEMEnOut275,MEMAddrOut275,MEMRWEnOut275
,MEMEnOut176,MEMDataOut76,MEMDataIn76,MEMAddrOut176,MEMRWEnOut176
,MEMEnOut276,MEMAddrOut276,MEMRWEnOut276
,MEMEnOut177,MEMDataOut77,MEMDataIn77,MEMAddrOut177,MEMRWEnOut177
,MEMEnOut277,MEMAddrOut277,MEMRWEnOut277
,MEMEnOut178,MEMDataOut78,MEMDataIn78,MEMAddrOut178,MEMRWEnOut178
,MEMEnOut278,MEMAddrOut278,MEMRWEnOut278
,MEMEnOut179,MEMDataOut79,MEMDataIn79,MEMAddrOut179,MEMRWEnOut179
,MEMEnOut279,MEMAddrOut279,MEMRWEnOut279
,MEMEnOut180,MEMDataOut80,MEMDataIn80,MEMAddrOut180,MEMRWEnOut180
,MEMEnOut280,MEMAddrOut280,MEMRWEnOut280
,MEMEnOut181,MEMDataOut81,MEMDataIn81,MEMAddrOut181,MEMRWEnOut181
,MEMEnOut281,MEMAddrOut281,MEMRWEnOut281
,MEMEnOut182,MEMDataOut82,MEMDataIn82,MEMAddrOut182,MEMRWEnOut182
,MEMEnOut282,MEMAddrOut282,MEMRWEnOut282
,MEMEnOut183,MEMDataOut83,MEMDataIn83,MEMAddrOut183,MEMRWEnOut183
,MEMEnOut283,MEMAddrOut283,MEMRWEnOut283
,MEMEnOut184,MEMDataOut84,MEMDataIn84,MEMAddrOut184,MEMRWEnOut184
,MEMEnOut284,MEMAddrOut284,MEMRWEnOut284
,MEMEnOut185,MEMDataOut85,MEMDataIn85,MEMAddrOut185,MEMRWEnOut185
,MEMEnOut285,MEMAddrOut285,MEMRWEnOut285
,MEMEnOut186,MEMDataOut86,MEMDataIn86,MEMAddrOut186,MEMRWEnOut186
,MEMEnOut286,MEMAddrOut286,MEMRWEnOut286
,MEMEnOut187,MEMDataOut87,MEMDataIn87,MEMAddrOut187,MEMRWEnOut187
,MEMEnOut287,MEMAddrOut287,MEMRWEnOut287
,MEMEnOut188,MEMDataOut88,MEMDataIn88,MEMAddrOut188,MEMRWEnOut188
,MEMEnOut288,MEMAddrOut288,MEMRWEnOut288
,MEMEnOut189,MEMDataOut89,MEMDataIn89,MEMAddrOut189,MEMRWEnOut189
,MEMEnOut289,MEMAddrOut289,MEMRWEnOut289
,MEMEnOut190,MEMDataOut90,MEMDataIn90,MEMAddrOut190,MEMRWEnOut190
,MEMEnOut290,MEMAddrOut290,MEMRWEnOut290
,MEMEnOut191,MEMDataOut91,MEMDataIn91,MEMAddrOut191,MEMRWEnOut191
,MEMEnOut291,MEMAddrOut291,MEMRWEnOut291
,MEMEnOut192,MEMDataOut92,MEMDataIn92,MEMAddrOut192,MEMRWEnOut192
,MEMEnOut292,MEMAddrOut292,MEMRWEnOut292
,MEMEnOut193,MEMDataOut93,MEMDataIn93,MEMAddrOut193,MEMRWEnOut193
,MEMEnOut293,MEMAddrOut293,MEMRWEnOut293
,MEMEnOut194,MEMDataOut94,MEMDataIn94,MEMAddrOut194,MEMRWEnOut194
,MEMEnOut294,MEMAddrOut294,MEMRWEnOut294
,MEMEnOut195,MEMDataOut95,MEMDataIn95,MEMAddrOut195,MEMRWEnOut195
,MEMEnOut295,MEMAddrOut295,MEMRWEnOut295
,MEMEnOut196,MEMDataOut96,MEMDataIn96,MEMAddrOut196,MEMRWEnOut196
,MEMEnOut296,MEMAddrOut296,MEMRWEnOut296
,MEMEnOut197,MEMDataOut97,MEMDataIn97,MEMAddrOut197,MEMRWEnOut197
,MEMEnOut297,MEMAddrOut297,MEMRWEnOut297
,MEMEnOut198,MEMDataOut98,MEMDataIn98,MEMAddrOut198,MEMRWEnOut198
,MEMEnOut298,MEMAddrOut298,MEMRWEnOut298
,MEMEnOut199,MEMDataOut99,MEMDataIn99,MEMAddrOut199,MEMRWEnOut199
,MEMEnOut299,MEMAddrOut299,MEMRWEnOut299
,MEMEnOut1100,MEMDataOut100,MEMDataIn100,MEMAddrOut1100,MEMRWEnOut1100
,MEMEnOut2100,MEMAddrOut2100,MEMRWEnOut2100
,MEMEnOut1101,MEMDataOut101,MEMDataIn101,MEMAddrOut1101,MEMRWEnOut1101
,MEMEnOut2101,MEMAddrOut2101,MEMRWEnOut2101
,MEMEnOut1102,MEMDataOut102,MEMDataIn102,MEMAddrOut1102,MEMRWEnOut1102
,MEMEnOut2102,MEMAddrOut2102,MEMRWEnOut2102
,MEMEnOut1103,MEMDataOut103,MEMDataIn103,MEMAddrOut1103,MEMRWEnOut1103
,MEMEnOut2103,MEMAddrOut2103,MEMRWEnOut2103
,MEMEnOut1104,MEMDataOut104,MEMDataIn104,MEMAddrOut1104,MEMRWEnOut1104
,MEMEnOut2104,MEMAddrOut2104,MEMRWEnOut2104
,MEMEnOut1105,MEMDataOut105,MEMDataIn105,MEMAddrOut1105,MEMRWEnOut1105
,MEMEnOut2105,MEMAddrOut2105,MEMRWEnOut2105
,MEMEnOut1106,MEMDataOut106,MEMDataIn106,MEMAddrOut1106,MEMRWEnOut1106
,MEMEnOut2106,MEMAddrOut2106,MEMRWEnOut2106
,MEMEnOut1107,MEMDataOut107,MEMDataIn107,MEMAddrOut1107,MEMRWEnOut1107
,MEMEnOut2107,MEMAddrOut2107,MEMRWEnOut2107);
input [3455:0] mLocalDataIn;
output [3455:0] mLocalDataOut;
input [38:0] mILocalDataIn;
output [38:0] mILocalDataOut;
input [107:0] MEMEnIn1;
input [107:0] MEMRWEnIn1;
input [647:0] MEMAddrIn1;
input IMEMEnIn1;
input IMEMRWEnIn1;
input [4:0] IMEMAddrIn1;
output IMEMEnOut1;
output IMEMRWEnOut1;
output [4:0] IMEMAddrOut1;
input [107:0] MEMEnIn2;
input [107:0] MEMRWEnIn2;
input [647:0] MEMAddrIn2;
input IMEMEnIn2;
input IMEMRWEnIn2;
input [4:0] IMEMAddrIn2;
output IMEMEnOut2;
output IMEMRWEnOut2;
output [4:0] IMEMAddrOut2;
output MEMEnOut10;
output MEMRWEnOut10;
output [31:0] MEMDataOut0;
input [31:0] MEMDataIn0;
output [5:0] MEMAddrOut10;
output MEMEnOut11;
output MEMRWEnOut11;
output [31:0] MEMDataOut1;
input [31:0] MEMDataIn1;
output [5:0] MEMAddrOut11;
output MEMEnOut12;
output MEMRWEnOut12;
output [31:0] MEMDataOut2;
input [31:0] MEMDataIn2;
output [5:0] MEMAddrOut12;
output MEMEnOut13;
output MEMRWEnOut13;
output [31:0] MEMDataOut3;
input [31:0] MEMDataIn3;
output [5:0] MEMAddrOut13;
output MEMEnOut14;
output MEMRWEnOut14;
output [31:0] MEMDataOut4;
input [31:0] MEMDataIn4;
output [5:0] MEMAddrOut14;
output MEMEnOut15;
output MEMRWEnOut15;
output [31:0] MEMDataOut5;
input [31:0] MEMDataIn5;
output [5:0] MEMAddrOut15;
output MEMEnOut16;
output MEMRWEnOut16;
output [31:0] MEMDataOut6;
input [31:0] MEMDataIn6;
output [5:0] MEMAddrOut16;
output MEMEnOut17;
output MEMRWEnOut17;
output [31:0] MEMDataOut7;
input [31:0] MEMDataIn7;
output [5:0] MEMAddrOut17;
output MEMEnOut18;
output MEMRWEnOut18;
output [31:0] MEMDataOut8;
input [31:0] MEMDataIn8;
output [5:0] MEMAddrOut18;
output MEMEnOut19;
output MEMRWEnOut19;
output [31:0] MEMDataOut9;
input [31:0] MEMDataIn9;
output [5:0] MEMAddrOut19;
output MEMEnOut110;
output MEMRWEnOut110;
output [31:0] MEMDataOut10;
input [31:0] MEMDataIn10;
output [5:0] MEMAddrOut110;
output MEMEnOut111;
output MEMRWEnOut111;
output [31:0] MEMDataOut11;
input [31:0] MEMDataIn11;
output [5:0] MEMAddrOut111;
output MEMEnOut112;
output MEMRWEnOut112;
output [31:0] MEMDataOut12;
input [31:0] MEMDataIn12;
output [5:0] MEMAddrOut112;
output MEMEnOut113;
output MEMRWEnOut113;
output [31:0] MEMDataOut13;
input [31:0] MEMDataIn13;
output [5:0] MEMAddrOut113;
output MEMEnOut114;
output MEMRWEnOut114;
output [31:0] MEMDataOut14;
input [31:0] MEMDataIn14;
output [5:0] MEMAddrOut114;
output MEMEnOut115;
output MEMRWEnOut115;
output [31:0] MEMDataOut15;
input [31:0] MEMDataIn15;
output [5:0] MEMAddrOut115;
output MEMEnOut116;
output MEMRWEnOut116;
output [31:0] MEMDataOut16;
input [31:0] MEMDataIn16;
output [5:0] MEMAddrOut116;
output MEMEnOut117;
output MEMRWEnOut117;
output [31:0] MEMDataOut17;
input [31:0] MEMDataIn17;
output [5:0] MEMAddrOut117;
output MEMEnOut118;
output MEMRWEnOut118;
output [31:0] MEMDataOut18;
input [31:0] MEMDataIn18;
output [5:0] MEMAddrOut118;
output MEMEnOut119;
output MEMRWEnOut119;
output [31:0] MEMDataOut19;
input [31:0] MEMDataIn19;
output [5:0] MEMAddrOut119;
output MEMEnOut120;
output MEMRWEnOut120;
output [31:0] MEMDataOut20;
input [31:0] MEMDataIn20;
output [5:0] MEMAddrOut120;
output MEMEnOut121;
output MEMRWEnOut121;
output [31:0] MEMDataOut21;
input [31:0] MEMDataIn21;
output [5:0] MEMAddrOut121;
output MEMEnOut122;
output MEMRWEnOut122;
output [31:0] MEMDataOut22;
input [31:0] MEMDataIn22;
output [5:0] MEMAddrOut122;
output MEMEnOut123;
output MEMRWEnOut123;
output [31:0] MEMDataOut23;
input [31:0] MEMDataIn23;
output [5:0] MEMAddrOut123;
output MEMEnOut124;
output MEMRWEnOut124;
output [31:0] MEMDataOut24;
input [31:0] MEMDataIn24;
output [5:0] MEMAddrOut124;
output MEMEnOut125;
output MEMRWEnOut125;
output [31:0] MEMDataOut25;
input [31:0] MEMDataIn25;
output [5:0] MEMAddrOut125;
output MEMEnOut126;
output MEMRWEnOut126;
output [31:0] MEMDataOut26;
input [31:0] MEMDataIn26;
output [5:0] MEMAddrOut126;
output MEMEnOut127;
output MEMRWEnOut127;
output [31:0] MEMDataOut27;
input [31:0] MEMDataIn27;
output [5:0] MEMAddrOut127;
output MEMEnOut128;
output MEMRWEnOut128;
output [31:0] MEMDataOut28;
input [31:0] MEMDataIn28;
output [5:0] MEMAddrOut128;
output MEMEnOut129;
output MEMRWEnOut129;
output [31:0] MEMDataOut29;
input [31:0] MEMDataIn29;
output [5:0] MEMAddrOut129;
output MEMEnOut130;
output MEMRWEnOut130;
output [31:0] MEMDataOut30;
input [31:0] MEMDataIn30;
output [5:0] MEMAddrOut130;
output MEMEnOut131;
output MEMRWEnOut131;
output [31:0] MEMDataOut31;
input [31:0] MEMDataIn31;
output [5:0] MEMAddrOut131;
output MEMEnOut132;
output MEMRWEnOut132;
output [31:0] MEMDataOut32;
input [31:0] MEMDataIn32;
output [5:0] MEMAddrOut132;
output MEMEnOut133;
output MEMRWEnOut133;
output [31:0] MEMDataOut33;
input [31:0] MEMDataIn33;
output [5:0] MEMAddrOut133;
output MEMEnOut134;
output MEMRWEnOut134;
output [31:0] MEMDataOut34;
input [31:0] MEMDataIn34;
output [5:0] MEMAddrOut134;
output MEMEnOut135;
output MEMRWEnOut135;
output [31:0] MEMDataOut35;
input [31:0] MEMDataIn35;
output [5:0] MEMAddrOut135;
output MEMEnOut136;
output MEMRWEnOut136;
output [31:0] MEMDataOut36;
input [31:0] MEMDataIn36;
output [5:0] MEMAddrOut136;
output MEMEnOut137;
output MEMRWEnOut137;
output [31:0] MEMDataOut37;
input [31:0] MEMDataIn37;
output [5:0] MEMAddrOut137;
output MEMEnOut138;
output MEMRWEnOut138;
output [31:0] MEMDataOut38;
input [31:0] MEMDataIn38;
output [5:0] MEMAddrOut138;
output MEMEnOut139;
output MEMRWEnOut139;
output [31:0] MEMDataOut39;
input [31:0] MEMDataIn39;
output [5:0] MEMAddrOut139;
output MEMEnOut140;
output MEMRWEnOut140;
output [31:0] MEMDataOut40;
input [31:0] MEMDataIn40;
output [5:0] MEMAddrOut140;
output MEMEnOut141;
output MEMRWEnOut141;
output [31:0] MEMDataOut41;
input [31:0] MEMDataIn41;
output [5:0] MEMAddrOut141;
output MEMEnOut142;
output MEMRWEnOut142;
output [31:0] MEMDataOut42;
input [31:0] MEMDataIn42;
output [5:0] MEMAddrOut142;
output MEMEnOut143;
output MEMRWEnOut143;
output [31:0] MEMDataOut43;
input [31:0] MEMDataIn43;
output [5:0] MEMAddrOut143;
output MEMEnOut144;
output MEMRWEnOut144;
output [31:0] MEMDataOut44;
input [31:0] MEMDataIn44;
output [5:0] MEMAddrOut144;
output MEMEnOut145;
output MEMRWEnOut145;
output [31:0] MEMDataOut45;
input [31:0] MEMDataIn45;
output [5:0] MEMAddrOut145;
output MEMEnOut146;
output MEMRWEnOut146;
output [31:0] MEMDataOut46;
input [31:0] MEMDataIn46;
output [5:0] MEMAddrOut146;
output MEMEnOut147;
output MEMRWEnOut147;
output [31:0] MEMDataOut47;
input [31:0] MEMDataIn47;
output [5:0] MEMAddrOut147;
output MEMEnOut148;
output MEMRWEnOut148;
output [31:0] MEMDataOut48;
input [31:0] MEMDataIn48;
output [5:0] MEMAddrOut148;
output MEMEnOut149;
output MEMRWEnOut149;
output [31:0] MEMDataOut49;
input [31:0] MEMDataIn49;
output [5:0] MEMAddrOut149;
output MEMEnOut150;
output MEMRWEnOut150;
output [31:0] MEMDataOut50;
input [31:0] MEMDataIn50;
output [5:0] MEMAddrOut150;
output MEMEnOut151;
output MEMRWEnOut151;
output [31:0] MEMDataOut51;
input [31:0] MEMDataIn51;
output [5:0] MEMAddrOut151;
output MEMEnOut152;
output MEMRWEnOut152;
output [31:0] MEMDataOut52;
input [31:0] MEMDataIn52;
output [5:0] MEMAddrOut152;
output MEMEnOut153;
output MEMRWEnOut153;
output [31:0] MEMDataOut53;
input [31:0] MEMDataIn53;
output [5:0] MEMAddrOut153;
output MEMEnOut154;
output MEMRWEnOut154;
output [31:0] MEMDataOut54;
input [31:0] MEMDataIn54;
output [5:0] MEMAddrOut154;
output MEMEnOut155;
output MEMRWEnOut155;
output [31:0] MEMDataOut55;
input [31:0] MEMDataIn55;
output [5:0] MEMAddrOut155;
output MEMEnOut156;
output MEMRWEnOut156;
output [31:0] MEMDataOut56;
input [31:0] MEMDataIn56;
output [5:0] MEMAddrOut156;
output MEMEnOut157;
output MEMRWEnOut157;
output [31:0] MEMDataOut57;
input [31:0] MEMDataIn57;
output [5:0] MEMAddrOut157;
output MEMEnOut158;
output MEMRWEnOut158;
output [31:0] MEMDataOut58;
input [31:0] MEMDataIn58;
output [5:0] MEMAddrOut158;
output MEMEnOut159;
output MEMRWEnOut159;
output [31:0] MEMDataOut59;
input [31:0] MEMDataIn59;
output [5:0] MEMAddrOut159;
output MEMEnOut160;
output MEMRWEnOut160;
output [31:0] MEMDataOut60;
input [31:0] MEMDataIn60;
output [5:0] MEMAddrOut160;
output MEMEnOut161;
output MEMRWEnOut161;
output [31:0] MEMDataOut61;
input [31:0] MEMDataIn61;
output [5:0] MEMAddrOut161;
output MEMEnOut162;
output MEMRWEnOut162;
output [31:0] MEMDataOut62;
input [31:0] MEMDataIn62;
output [5:0] MEMAddrOut162;
output MEMEnOut163;
output MEMRWEnOut163;
output [31:0] MEMDataOut63;
input [31:0] MEMDataIn63;
output [5:0] MEMAddrOut163;
output MEMEnOut164;
output MEMRWEnOut164;
output [31:0] MEMDataOut64;
input [31:0] MEMDataIn64;
output [5:0] MEMAddrOut164;
output MEMEnOut165;
output MEMRWEnOut165;
output [31:0] MEMDataOut65;
input [31:0] MEMDataIn65;
output [5:0] MEMAddrOut165;
output MEMEnOut166;
output MEMRWEnOut166;
output [31:0] MEMDataOut66;
input [31:0] MEMDataIn66;
output [5:0] MEMAddrOut166;
output MEMEnOut167;
output MEMRWEnOut167;
output [31:0] MEMDataOut67;
input [31:0] MEMDataIn67;
output [5:0] MEMAddrOut167;
output MEMEnOut168;
output MEMRWEnOut168;
output [31:0] MEMDataOut68;
input [31:0] MEMDataIn68;
output [5:0] MEMAddrOut168;
output MEMEnOut169;
output MEMRWEnOut169;
output [31:0] MEMDataOut69;
input [31:0] MEMDataIn69;
output [5:0] MEMAddrOut169;
output MEMEnOut170;
output MEMRWEnOut170;
output [31:0] MEMDataOut70;
input [31:0] MEMDataIn70;
output [5:0] MEMAddrOut170;
output MEMEnOut171;
output MEMRWEnOut171;
output [31:0] MEMDataOut71;
input [31:0] MEMDataIn71;
output [5:0] MEMAddrOut171;
output MEMEnOut172;
output MEMRWEnOut172;
output [31:0] MEMDataOut72;
input [31:0] MEMDataIn72;
output [5:0] MEMAddrOut172;
output MEMEnOut173;
output MEMRWEnOut173;
output [31:0] MEMDataOut73;
input [31:0] MEMDataIn73;
output [5:0] MEMAddrOut173;
output MEMEnOut174;
output MEMRWEnOut174;
output [31:0] MEMDataOut74;
input [31:0] MEMDataIn74;
output [5:0] MEMAddrOut174;
output MEMEnOut175;
output MEMRWEnOut175;
output [31:0] MEMDataOut75;
input [31:0] MEMDataIn75;
output [5:0] MEMAddrOut175;
output MEMEnOut176;
output MEMRWEnOut176;
output [31:0] MEMDataOut76;
input [31:0] MEMDataIn76;
output [5:0] MEMAddrOut176;
output MEMEnOut177;
output MEMRWEnOut177;
output [31:0] MEMDataOut77;
input [31:0] MEMDataIn77;
output [5:0] MEMAddrOut177;
output MEMEnOut178;
output MEMRWEnOut178;
output [31:0] MEMDataOut78;
input [31:0] MEMDataIn78;
output [5:0] MEMAddrOut178;
output MEMEnOut179;
output MEMRWEnOut179;
output [31:0] MEMDataOut79;
input [31:0] MEMDataIn79;
output [5:0] MEMAddrOut179;
output MEMEnOut180;
output MEMRWEnOut180;
output [31:0] MEMDataOut80;
input [31:0] MEMDataIn80;
output [5:0] MEMAddrOut180;
output MEMEnOut181;
output MEMRWEnOut181;
output [31:0] MEMDataOut81;
input [31:0] MEMDataIn81;
output [5:0] MEMAddrOut181;
output MEMEnOut182;
output MEMRWEnOut182;
output [31:0] MEMDataOut82;
input [31:0] MEMDataIn82;
output [5:0] MEMAddrOut182;
output MEMEnOut183;
output MEMRWEnOut183;
output [31:0] MEMDataOut83;
input [31:0] MEMDataIn83;
output [5:0] MEMAddrOut183;
output MEMEnOut184;
output MEMRWEnOut184;
output [31:0] MEMDataOut84;
input [31:0] MEMDataIn84;
output [5:0] MEMAddrOut184;
output MEMEnOut185;
output MEMRWEnOut185;
output [31:0] MEMDataOut85;
input [31:0] MEMDataIn85;
output [5:0] MEMAddrOut185;
output MEMEnOut186;
output MEMRWEnOut186;
output [31:0] MEMDataOut86;
input [31:0] MEMDataIn86;
output [5:0] MEMAddrOut186;
output MEMEnOut187;
output MEMRWEnOut187;
output [31:0] MEMDataOut87;
input [31:0] MEMDataIn87;
output [5:0] MEMAddrOut187;
output MEMEnOut188;
output MEMRWEnOut188;
output [31:0] MEMDataOut88;
input [31:0] MEMDataIn88;
output [5:0] MEMAddrOut188;
output MEMEnOut189;
output MEMRWEnOut189;
output [31:0] MEMDataOut89;
input [31:0] MEMDataIn89;
output [5:0] MEMAddrOut189;
output MEMEnOut190;
output MEMRWEnOut190;
output [31:0] MEMDataOut90;
input [31:0] MEMDataIn90;
output [5:0] MEMAddrOut190;
output MEMEnOut191;
output MEMRWEnOut191;
output [31:0] MEMDataOut91;
input [31:0] MEMDataIn91;
output [5:0] MEMAddrOut191;
output MEMEnOut192;
output MEMRWEnOut192;
output [31:0] MEMDataOut92;
input [31:0] MEMDataIn92;
output [5:0] MEMAddrOut192;
output MEMEnOut193;
output MEMRWEnOut193;
output [31:0] MEMDataOut93;
input [31:0] MEMDataIn93;
output [5:0] MEMAddrOut193;
output MEMEnOut194;
output MEMRWEnOut194;
output [31:0] MEMDataOut94;
input [31:0] MEMDataIn94;
output [5:0] MEMAddrOut194;
output MEMEnOut195;
output MEMRWEnOut195;
output [31:0] MEMDataOut95;
input [31:0] MEMDataIn95;
output [5:0] MEMAddrOut195;
output MEMEnOut196;
output MEMRWEnOut196;
output [31:0] MEMDataOut96;
input [31:0] MEMDataIn96;
output [5:0] MEMAddrOut196;
output MEMEnOut197;
output MEMRWEnOut197;
output [31:0] MEMDataOut97;
input [31:0] MEMDataIn97;
output [5:0] MEMAddrOut197;
output MEMEnOut198;
output MEMRWEnOut198;
output [31:0] MEMDataOut98;
input [31:0] MEMDataIn98;
output [5:0] MEMAddrOut198;
output MEMEnOut199;
output MEMRWEnOut199;
output [31:0] MEMDataOut99;
input [31:0] MEMDataIn99;
output [5:0] MEMAddrOut199;
output MEMEnOut1100;
output MEMRWEnOut1100;
output [31:0] MEMDataOut100;
input [31:0] MEMDataIn100;
output [5:0] MEMAddrOut1100;
output MEMEnOut1101;
output MEMRWEnOut1101;
output [31:0] MEMDataOut101;
input [31:0] MEMDataIn101;
output [5:0] MEMAddrOut1101;
output MEMEnOut1102;
output MEMRWEnOut1102;
output [31:0] MEMDataOut102;
input [31:0] MEMDataIn102;
output [5:0] MEMAddrOut1102;
output MEMEnOut1103;
output MEMRWEnOut1103;
output [31:0] MEMDataOut103;
input [31:0] MEMDataIn103;
output [5:0] MEMAddrOut1103;
output MEMEnOut1104;
output MEMRWEnOut1104;
output [31:0] MEMDataOut104;
input [31:0] MEMDataIn104;
output [5:0] MEMAddrOut1104;
output MEMEnOut1105;
output MEMRWEnOut1105;
output [31:0] MEMDataOut105;
input [31:0] MEMDataIn105;
output [5:0] MEMAddrOut1105;
output MEMEnOut1106;
output MEMRWEnOut1106;
output [31:0] MEMDataOut106;
input [31:0] MEMDataIn106;
output [5:0] MEMAddrOut1106;
output MEMEnOut1107;
output MEMRWEnOut1107;
output [31:0] MEMDataOut107;
input [31:0] MEMDataIn107;
output [5:0] MEMAddrOut1107;
assign MEMEnOut10= MEMEnIn1[0:0];
assign MEMRWEnOut10= MEMRWEnIn1[0:0];
assign MEMDataOut0= mLocalDataIn[31:0];
assign mLocalDataOut[31:0] = MEMDataIn0;
assign MEMAddrOut10= MEMAddrIn1[5:0];
assign MEMEnOut11= MEMEnIn1[1:1];
assign MEMRWEnOut11= MEMRWEnIn1[1:1];
assign MEMDataOut1= mLocalDataIn[63:32];
assign mLocalDataOut[63:32] = MEMDataIn1;
assign MEMAddrOut11= MEMAddrIn1[11:6];
assign MEMEnOut12= MEMEnIn1[2:2];
assign MEMRWEnOut12= MEMRWEnIn1[2:2];
assign MEMDataOut2= mLocalDataIn[95:64];
assign mLocalDataOut[95:64] = MEMDataIn2;
assign MEMAddrOut12= MEMAddrIn1[17:12];
assign MEMEnOut13= MEMEnIn1[3:3];
assign MEMRWEnOut13= MEMRWEnIn1[3:3];
assign MEMDataOut3= mLocalDataIn[127:96];
assign mLocalDataOut[127:96] = MEMDataIn3;
assign MEMAddrOut13= MEMAddrIn1[23:18];
assign MEMEnOut14= MEMEnIn1[4:4];
assign MEMRWEnOut14= MEMRWEnIn1[4:4];
assign MEMDataOut4= mLocalDataIn[159:128];
assign mLocalDataOut[159:128] = MEMDataIn4;
assign MEMAddrOut14= MEMAddrIn1[29:24];
assign MEMEnOut15= MEMEnIn1[5:5];
assign MEMRWEnOut15= MEMRWEnIn1[5:5];
assign MEMDataOut5= mLocalDataIn[191:160];
assign mLocalDataOut[191:160] = MEMDataIn5;
assign MEMAddrOut15= MEMAddrIn1[35:30];
assign MEMEnOut16= MEMEnIn1[6:6];
assign MEMRWEnOut16= MEMRWEnIn1[6:6];
assign MEMDataOut6= mLocalDataIn[223:192];
assign mLocalDataOut[223:192] = MEMDataIn6;
assign MEMAddrOut16= MEMAddrIn1[41:36];
assign MEMEnOut17= MEMEnIn1[7:7];
assign MEMRWEnOut17= MEMRWEnIn1[7:7];
assign MEMDataOut7= mLocalDataIn[255:224];
assign mLocalDataOut[255:224] = MEMDataIn7;
assign MEMAddrOut17= MEMAddrIn1[47:42];
assign MEMEnOut18= MEMEnIn1[8:8];
assign MEMRWEnOut18= MEMRWEnIn1[8:8];
assign MEMDataOut8= mLocalDataIn[287:256];
assign mLocalDataOut[287:256] = MEMDataIn8;
assign MEMAddrOut18= MEMAddrIn1[53:48];
assign MEMEnOut19= MEMEnIn1[9:9];
assign MEMRWEnOut19= MEMRWEnIn1[9:9];
assign MEMDataOut9= mLocalDataIn[319:288];
assign mLocalDataOut[319:288] = MEMDataIn9;
assign MEMAddrOut19= MEMAddrIn1[59:54];
assign MEMEnOut110= MEMEnIn1[10:10];
assign MEMRWEnOut110= MEMRWEnIn1[10:10];
assign MEMDataOut10= mLocalDataIn[351:320];
assign mLocalDataOut[351:320] = MEMDataIn10;
assign MEMAddrOut110= MEMAddrIn1[65:60];
assign MEMEnOut111= MEMEnIn1[11:11];
assign MEMRWEnOut111= MEMRWEnIn1[11:11];
assign MEMDataOut11= mLocalDataIn[383:352];
assign mLocalDataOut[383:352] = MEMDataIn11;
assign MEMAddrOut111= MEMAddrIn1[71:66];
assign MEMEnOut112= MEMEnIn1[12:12];
assign MEMRWEnOut112= MEMRWEnIn1[12:12];
assign MEMDataOut12= mLocalDataIn[415:384];
assign mLocalDataOut[415:384] = MEMDataIn12;
assign MEMAddrOut112= MEMAddrIn1[77:72];
assign MEMEnOut113= MEMEnIn1[13:13];
assign MEMRWEnOut113= MEMRWEnIn1[13:13];
assign MEMDataOut13= mLocalDataIn[447:416];
assign mLocalDataOut[447:416] = MEMDataIn13;
assign MEMAddrOut113= MEMAddrIn1[83:78];
assign MEMEnOut114= MEMEnIn1[14:14];
assign MEMRWEnOut114= MEMRWEnIn1[14:14];
assign MEMDataOut14= mLocalDataIn[479:448];
assign mLocalDataOut[479:448] = MEMDataIn14;
assign MEMAddrOut114= MEMAddrIn1[89:84];
assign MEMEnOut115= MEMEnIn1[15:15];
assign MEMRWEnOut115= MEMRWEnIn1[15:15];
assign MEMDataOut15= mLocalDataIn[511:480];
assign mLocalDataOut[511:480] = MEMDataIn15;
assign MEMAddrOut115= MEMAddrIn1[95:90];
assign MEMEnOut116= MEMEnIn1[16:16];
assign MEMRWEnOut116= MEMRWEnIn1[16:16];
assign MEMDataOut16= mLocalDataIn[543:512];
assign mLocalDataOut[543:512] = MEMDataIn16;
assign MEMAddrOut116= MEMAddrIn1[101:96];
assign MEMEnOut117= MEMEnIn1[17:17];
assign MEMRWEnOut117= MEMRWEnIn1[17:17];
assign MEMDataOut17= mLocalDataIn[575:544];
assign mLocalDataOut[575:544] = MEMDataIn17;
assign MEMAddrOut117= MEMAddrIn1[107:102];
assign MEMEnOut118= MEMEnIn1[18:18];
assign MEMRWEnOut118= MEMRWEnIn1[18:18];
assign MEMDataOut18= mLocalDataIn[607:576];
assign mLocalDataOut[607:576] = MEMDataIn18;
assign MEMAddrOut118= MEMAddrIn1[113:108];
assign MEMEnOut119= MEMEnIn1[19:19];
assign MEMRWEnOut119= MEMRWEnIn1[19:19];
assign MEMDataOut19= mLocalDataIn[639:608];
assign mLocalDataOut[639:608] = MEMDataIn19;
assign MEMAddrOut119= MEMAddrIn1[119:114];
assign MEMEnOut120= MEMEnIn1[20:20];
assign MEMRWEnOut120= MEMRWEnIn1[20:20];
assign MEMDataOut20= mLocalDataIn[671:640];
assign mLocalDataOut[671:640] = MEMDataIn20;
assign MEMAddrOut120= MEMAddrIn1[125:120];
assign MEMEnOut121= MEMEnIn1[21:21];
assign MEMRWEnOut121= MEMRWEnIn1[21:21];
assign MEMDataOut21= mLocalDataIn[703:672];
assign mLocalDataOut[703:672] = MEMDataIn21;
assign MEMAddrOut121= MEMAddrIn1[131:126];
assign MEMEnOut122= MEMEnIn1[22:22];
assign MEMRWEnOut122= MEMRWEnIn1[22:22];
assign MEMDataOut22= mLocalDataIn[735:704];
assign mLocalDataOut[735:704] = MEMDataIn22;
assign MEMAddrOut122= MEMAddrIn1[137:132];
assign MEMEnOut123= MEMEnIn1[23:23];
assign MEMRWEnOut123= MEMRWEnIn1[23:23];
assign MEMDataOut23= mLocalDataIn[767:736];
assign mLocalDataOut[767:736] = MEMDataIn23;
assign MEMAddrOut123= MEMAddrIn1[143:138];
assign MEMEnOut124= MEMEnIn1[24:24];
assign MEMRWEnOut124= MEMRWEnIn1[24:24];
assign MEMDataOut24= mLocalDataIn[799:768];
assign mLocalDataOut[799:768] = MEMDataIn24;
assign MEMAddrOut124= MEMAddrIn1[149:144];
assign MEMEnOut125= MEMEnIn1[25:25];
assign MEMRWEnOut125= MEMRWEnIn1[25:25];
assign MEMDataOut25= mLocalDataIn[831:800];
assign mLocalDataOut[831:800] = MEMDataIn25;
assign MEMAddrOut125= MEMAddrIn1[155:150];
assign MEMEnOut126= MEMEnIn1[26:26];
assign MEMRWEnOut126= MEMRWEnIn1[26:26];
assign MEMDataOut26= mLocalDataIn[863:832];
assign mLocalDataOut[863:832] = MEMDataIn26;
assign MEMAddrOut126= MEMAddrIn1[161:156];
assign MEMEnOut127= MEMEnIn1[27:27];
assign MEMRWEnOut127= MEMRWEnIn1[27:27];
assign MEMDataOut27= mLocalDataIn[895:864];
assign mLocalDataOut[895:864] = MEMDataIn27;
assign MEMAddrOut127= MEMAddrIn1[167:162];
assign MEMEnOut128= MEMEnIn1[28:28];
assign MEMRWEnOut128= MEMRWEnIn1[28:28];
assign MEMDataOut28= mLocalDataIn[927:896];
assign mLocalDataOut[927:896] = MEMDataIn28;
assign MEMAddrOut128= MEMAddrIn1[173:168];
assign MEMEnOut129= MEMEnIn1[29:29];
assign MEMRWEnOut129= MEMRWEnIn1[29:29];
assign MEMDataOut29= mLocalDataIn[959:928];
assign mLocalDataOut[959:928] = MEMDataIn29;
assign MEMAddrOut129= MEMAddrIn1[179:174];
assign MEMEnOut130= MEMEnIn1[30:30];
assign MEMRWEnOut130= MEMRWEnIn1[30:30];
assign MEMDataOut30= mLocalDataIn[991:960];
assign mLocalDataOut[991:960] = MEMDataIn30;
assign MEMAddrOut130= MEMAddrIn1[185:180];
assign MEMEnOut131= MEMEnIn1[31:31];
assign MEMRWEnOut131= MEMRWEnIn1[31:31];
assign MEMDataOut31= mLocalDataIn[1023:992];
assign mLocalDataOut[1023:992] = MEMDataIn31;
assign MEMAddrOut131= MEMAddrIn1[191:186];
assign MEMEnOut132= MEMEnIn1[32:32];
assign MEMRWEnOut132= MEMRWEnIn1[32:32];
assign MEMDataOut32= mLocalDataIn[1055:1024];
assign mLocalDataOut[1055:1024] = MEMDataIn32;
assign MEMAddrOut132= MEMAddrIn1[197:192];
assign MEMEnOut133= MEMEnIn1[33:33];
assign MEMRWEnOut133= MEMRWEnIn1[33:33];
assign MEMDataOut33= mLocalDataIn[1087:1056];
assign mLocalDataOut[1087:1056] = MEMDataIn33;
assign MEMAddrOut133= MEMAddrIn1[203:198];
assign MEMEnOut134= MEMEnIn1[34:34];
assign MEMRWEnOut134= MEMRWEnIn1[34:34];
assign MEMDataOut34= mLocalDataIn[1119:1088];
assign mLocalDataOut[1119:1088] = MEMDataIn34;
assign MEMAddrOut134= MEMAddrIn1[209:204];
assign MEMEnOut135= MEMEnIn1[35:35];
assign MEMRWEnOut135= MEMRWEnIn1[35:35];
assign MEMDataOut35= mLocalDataIn[1151:1120];
assign mLocalDataOut[1151:1120] = MEMDataIn35;
assign MEMAddrOut135= MEMAddrIn1[215:210];
assign MEMEnOut136= MEMEnIn1[36:36];
assign MEMRWEnOut136= MEMRWEnIn1[36:36];
assign MEMDataOut36= mLocalDataIn[1183:1152];
assign mLocalDataOut[1183:1152] = MEMDataIn36;
assign MEMAddrOut136= MEMAddrIn1[221:216];
assign MEMEnOut137= MEMEnIn1[37:37];
assign MEMRWEnOut137= MEMRWEnIn1[37:37];
assign MEMDataOut37= mLocalDataIn[1215:1184];
assign mLocalDataOut[1215:1184] = MEMDataIn37;
assign MEMAddrOut137= MEMAddrIn1[227:222];
assign MEMEnOut138= MEMEnIn1[38:38];
assign MEMRWEnOut138= MEMRWEnIn1[38:38];
assign MEMDataOut38= mLocalDataIn[1247:1216];
assign mLocalDataOut[1247:1216] = MEMDataIn38;
assign MEMAddrOut138= MEMAddrIn1[233:228];
assign MEMEnOut139= MEMEnIn1[39:39];
assign MEMRWEnOut139= MEMRWEnIn1[39:39];
assign MEMDataOut39= mLocalDataIn[1279:1248];
assign mLocalDataOut[1279:1248] = MEMDataIn39;
assign MEMAddrOut139= MEMAddrIn1[239:234];
assign MEMEnOut140= MEMEnIn1[40:40];
assign MEMRWEnOut140= MEMRWEnIn1[40:40];
assign MEMDataOut40= mLocalDataIn[1311:1280];
assign mLocalDataOut[1311:1280] = MEMDataIn40;
assign MEMAddrOut140= MEMAddrIn1[245:240];
assign MEMEnOut141= MEMEnIn1[41:41];
assign MEMRWEnOut141= MEMRWEnIn1[41:41];
assign MEMDataOut41= mLocalDataIn[1343:1312];
assign mLocalDataOut[1343:1312] = MEMDataIn41;
assign MEMAddrOut141= MEMAddrIn1[251:246];
assign MEMEnOut142= MEMEnIn1[42:42];
assign MEMRWEnOut142= MEMRWEnIn1[42:42];
assign MEMDataOut42= mLocalDataIn[1375:1344];
assign mLocalDataOut[1375:1344] = MEMDataIn42;
assign MEMAddrOut142= MEMAddrIn1[257:252];
assign MEMEnOut143= MEMEnIn1[43:43];
assign MEMRWEnOut143= MEMRWEnIn1[43:43];
assign MEMDataOut43= mLocalDataIn[1407:1376];
assign mLocalDataOut[1407:1376] = MEMDataIn43;
assign MEMAddrOut143= MEMAddrIn1[263:258];
assign MEMEnOut144= MEMEnIn1[44:44];
assign MEMRWEnOut144= MEMRWEnIn1[44:44];
assign MEMDataOut44= mLocalDataIn[1439:1408];
assign mLocalDataOut[1439:1408] = MEMDataIn44;
assign MEMAddrOut144= MEMAddrIn1[269:264];
assign MEMEnOut145= MEMEnIn1[45:45];
assign MEMRWEnOut145= MEMRWEnIn1[45:45];
assign MEMDataOut45= mLocalDataIn[1471:1440];
assign mLocalDataOut[1471:1440] = MEMDataIn45;
assign MEMAddrOut145= MEMAddrIn1[275:270];
assign MEMEnOut146= MEMEnIn1[46:46];
assign MEMRWEnOut146= MEMRWEnIn1[46:46];
assign MEMDataOut46= mLocalDataIn[1503:1472];
assign mLocalDataOut[1503:1472] = MEMDataIn46;
assign MEMAddrOut146= MEMAddrIn1[281:276];
assign MEMEnOut147= MEMEnIn1[47:47];
assign MEMRWEnOut147= MEMRWEnIn1[47:47];
assign MEMDataOut47= mLocalDataIn[1535:1504];
assign mLocalDataOut[1535:1504] = MEMDataIn47;
assign MEMAddrOut147= MEMAddrIn1[287:282];
assign MEMEnOut148= MEMEnIn1[48:48];
assign MEMRWEnOut148= MEMRWEnIn1[48:48];
assign MEMDataOut48= mLocalDataIn[1567:1536];
assign mLocalDataOut[1567:1536] = MEMDataIn48;
assign MEMAddrOut148= MEMAddrIn1[293:288];
assign MEMEnOut149= MEMEnIn1[49:49];
assign MEMRWEnOut149= MEMRWEnIn1[49:49];
assign MEMDataOut49= mLocalDataIn[1599:1568];
assign mLocalDataOut[1599:1568] = MEMDataIn49;
assign MEMAddrOut149= MEMAddrIn1[299:294];
assign MEMEnOut150= MEMEnIn1[50:50];
assign MEMRWEnOut150= MEMRWEnIn1[50:50];
assign MEMDataOut50= mLocalDataIn[1631:1600];
assign mLocalDataOut[1631:1600] = MEMDataIn50;
assign MEMAddrOut150= MEMAddrIn1[305:300];
assign MEMEnOut151= MEMEnIn1[51:51];
assign MEMRWEnOut151= MEMRWEnIn1[51:51];
assign MEMDataOut51= mLocalDataIn[1663:1632];
assign mLocalDataOut[1663:1632] = MEMDataIn51;
assign MEMAddrOut151= MEMAddrIn1[311:306];
assign MEMEnOut152= MEMEnIn1[52:52];
assign MEMRWEnOut152= MEMRWEnIn1[52:52];
assign MEMDataOut52= mLocalDataIn[1695:1664];
assign mLocalDataOut[1695:1664] = MEMDataIn52;
assign MEMAddrOut152= MEMAddrIn1[317:312];
assign MEMEnOut153= MEMEnIn1[53:53];
assign MEMRWEnOut153= MEMRWEnIn1[53:53];
assign MEMDataOut53= mLocalDataIn[1727:1696];
assign mLocalDataOut[1727:1696] = MEMDataIn53;
assign MEMAddrOut153= MEMAddrIn1[323:318];
assign MEMEnOut154= MEMEnIn1[54:54];
assign MEMRWEnOut154= MEMRWEnIn1[54:54];
assign MEMDataOut54= mLocalDataIn[1759:1728];
assign mLocalDataOut[1759:1728] = MEMDataIn54;
assign MEMAddrOut154= MEMAddrIn1[329:324];
assign MEMEnOut155= MEMEnIn1[55:55];
assign MEMRWEnOut155= MEMRWEnIn1[55:55];
assign MEMDataOut55= mLocalDataIn[1791:1760];
assign mLocalDataOut[1791:1760] = MEMDataIn55;
assign MEMAddrOut155= MEMAddrIn1[335:330];
assign MEMEnOut156= MEMEnIn1[56:56];
assign MEMRWEnOut156= MEMRWEnIn1[56:56];
assign MEMDataOut56= mLocalDataIn[1823:1792];
assign mLocalDataOut[1823:1792] = MEMDataIn56;
assign MEMAddrOut156= MEMAddrIn1[341:336];
assign MEMEnOut157= MEMEnIn1[57:57];
assign MEMRWEnOut157= MEMRWEnIn1[57:57];
assign MEMDataOut57= mLocalDataIn[1855:1824];
assign mLocalDataOut[1855:1824] = MEMDataIn57;
assign MEMAddrOut157= MEMAddrIn1[347:342];
assign MEMEnOut158= MEMEnIn1[58:58];
assign MEMRWEnOut158= MEMRWEnIn1[58:58];
assign MEMDataOut58= mLocalDataIn[1887:1856];
assign mLocalDataOut[1887:1856] = MEMDataIn58;
assign MEMAddrOut158= MEMAddrIn1[353:348];
assign MEMEnOut159= MEMEnIn1[59:59];
assign MEMRWEnOut159= MEMRWEnIn1[59:59];
assign MEMDataOut59= mLocalDataIn[1919:1888];
assign mLocalDataOut[1919:1888] = MEMDataIn59;
assign MEMAddrOut159= MEMAddrIn1[359:354];
assign MEMEnOut160= MEMEnIn1[60:60];
assign MEMRWEnOut160= MEMRWEnIn1[60:60];
assign MEMDataOut60= mLocalDataIn[1951:1920];
assign mLocalDataOut[1951:1920] = MEMDataIn60;
assign MEMAddrOut160= MEMAddrIn1[365:360];
assign MEMEnOut161= MEMEnIn1[61:61];
assign MEMRWEnOut161= MEMRWEnIn1[61:61];
assign MEMDataOut61= mLocalDataIn[1983:1952];
assign mLocalDataOut[1983:1952] = MEMDataIn61;
assign MEMAddrOut161= MEMAddrIn1[371:366];
assign MEMEnOut162= MEMEnIn1[62:62];
assign MEMRWEnOut162= MEMRWEnIn1[62:62];
assign MEMDataOut62= mLocalDataIn[2015:1984];
assign mLocalDataOut[2015:1984] = MEMDataIn62;
assign MEMAddrOut162= MEMAddrIn1[377:372];
assign MEMEnOut163= MEMEnIn1[63:63];
assign MEMRWEnOut163= MEMRWEnIn1[63:63];
assign MEMDataOut63= mLocalDataIn[2047:2016];
assign mLocalDataOut[2047:2016] = MEMDataIn63;
assign MEMAddrOut163= MEMAddrIn1[383:378];
assign MEMEnOut164= MEMEnIn1[64:64];
assign MEMRWEnOut164= MEMRWEnIn1[64:64];
assign MEMDataOut64= mLocalDataIn[2079:2048];
assign mLocalDataOut[2079:2048] = MEMDataIn64;
assign MEMAddrOut164= MEMAddrIn1[389:384];
assign MEMEnOut165= MEMEnIn1[65:65];
assign MEMRWEnOut165= MEMRWEnIn1[65:65];
assign MEMDataOut65= mLocalDataIn[2111:2080];
assign mLocalDataOut[2111:2080] = MEMDataIn65;
assign MEMAddrOut165= MEMAddrIn1[395:390];
assign MEMEnOut166= MEMEnIn1[66:66];
assign MEMRWEnOut166= MEMRWEnIn1[66:66];
assign MEMDataOut66= mLocalDataIn[2143:2112];
assign mLocalDataOut[2143:2112] = MEMDataIn66;
assign MEMAddrOut166= MEMAddrIn1[401:396];
assign MEMEnOut167= MEMEnIn1[67:67];
assign MEMRWEnOut167= MEMRWEnIn1[67:67];
assign MEMDataOut67= mLocalDataIn[2175:2144];
assign mLocalDataOut[2175:2144] = MEMDataIn67;
assign MEMAddrOut167= MEMAddrIn1[407:402];
assign MEMEnOut168= MEMEnIn1[68:68];
assign MEMRWEnOut168= MEMRWEnIn1[68:68];
assign MEMDataOut68= mLocalDataIn[2207:2176];
assign mLocalDataOut[2207:2176] = MEMDataIn68;
assign MEMAddrOut168= MEMAddrIn1[413:408];
assign MEMEnOut169= MEMEnIn1[69:69];
assign MEMRWEnOut169= MEMRWEnIn1[69:69];
assign MEMDataOut69= mLocalDataIn[2239:2208];
assign mLocalDataOut[2239:2208] = MEMDataIn69;
assign MEMAddrOut169= MEMAddrIn1[419:414];
assign MEMEnOut170= MEMEnIn1[70:70];
assign MEMRWEnOut170= MEMRWEnIn1[70:70];
assign MEMDataOut70= mLocalDataIn[2271:2240];
assign mLocalDataOut[2271:2240] = MEMDataIn70;
assign MEMAddrOut170= MEMAddrIn1[425:420];
assign MEMEnOut171= MEMEnIn1[71:71];
assign MEMRWEnOut171= MEMRWEnIn1[71:71];
assign MEMDataOut71= mLocalDataIn[2303:2272];
assign mLocalDataOut[2303:2272] = MEMDataIn71;
assign MEMAddrOut171= MEMAddrIn1[431:426];
assign MEMEnOut172= MEMEnIn1[72:72];
assign MEMRWEnOut172= MEMRWEnIn1[72:72];
assign MEMDataOut72= mLocalDataIn[2335:2304];
assign mLocalDataOut[2335:2304] = MEMDataIn72;
assign MEMAddrOut172= MEMAddrIn1[437:432];
assign MEMEnOut173= MEMEnIn1[73:73];
assign MEMRWEnOut173= MEMRWEnIn1[73:73];
assign MEMDataOut73= mLocalDataIn[2367:2336];
assign mLocalDataOut[2367:2336] = MEMDataIn73;
assign MEMAddrOut173= MEMAddrIn1[443:438];
assign MEMEnOut174= MEMEnIn1[74:74];
assign MEMRWEnOut174= MEMRWEnIn1[74:74];
assign MEMDataOut74= mLocalDataIn[2399:2368];
assign mLocalDataOut[2399:2368] = MEMDataIn74;
assign MEMAddrOut174= MEMAddrIn1[449:444];
assign MEMEnOut175= MEMEnIn1[75:75];
assign MEMRWEnOut175= MEMRWEnIn1[75:75];
assign MEMDataOut75= mLocalDataIn[2431:2400];
assign mLocalDataOut[2431:2400] = MEMDataIn75;
assign MEMAddrOut175= MEMAddrIn1[455:450];
assign MEMEnOut176= MEMEnIn1[76:76];
assign MEMRWEnOut176= MEMRWEnIn1[76:76];
assign MEMDataOut76= mLocalDataIn[2463:2432];
assign mLocalDataOut[2463:2432] = MEMDataIn76;
assign MEMAddrOut176= MEMAddrIn1[461:456];
assign MEMEnOut177= MEMEnIn1[77:77];
assign MEMRWEnOut177= MEMRWEnIn1[77:77];
assign MEMDataOut77= mLocalDataIn[2495:2464];
assign mLocalDataOut[2495:2464] = MEMDataIn77;
assign MEMAddrOut177= MEMAddrIn1[467:462];
assign MEMEnOut178= MEMEnIn1[78:78];
assign MEMRWEnOut178= MEMRWEnIn1[78:78];
assign MEMDataOut78= mLocalDataIn[2527:2496];
assign mLocalDataOut[2527:2496] = MEMDataIn78;
assign MEMAddrOut178= MEMAddrIn1[473:468];
assign MEMEnOut179= MEMEnIn1[79:79];
assign MEMRWEnOut179= MEMRWEnIn1[79:79];
assign MEMDataOut79= mLocalDataIn[2559:2528];
assign mLocalDataOut[2559:2528] = MEMDataIn79;
assign MEMAddrOut179= MEMAddrIn1[479:474];
assign MEMEnOut180= MEMEnIn1[80:80];
assign MEMRWEnOut180= MEMRWEnIn1[80:80];
assign MEMDataOut80= mLocalDataIn[2591:2560];
assign mLocalDataOut[2591:2560] = MEMDataIn80;
assign MEMAddrOut180= MEMAddrIn1[485:480];
assign MEMEnOut181= MEMEnIn1[81:81];
assign MEMRWEnOut181= MEMRWEnIn1[81:81];
assign MEMDataOut81= mLocalDataIn[2623:2592];
assign mLocalDataOut[2623:2592] = MEMDataIn81;
assign MEMAddrOut181= MEMAddrIn1[491:486];
assign MEMEnOut182= MEMEnIn1[82:82];
assign MEMRWEnOut182= MEMRWEnIn1[82:82];
assign MEMDataOut82= mLocalDataIn[2655:2624];
assign mLocalDataOut[2655:2624] = MEMDataIn82;
assign MEMAddrOut182= MEMAddrIn1[497:492];
assign MEMEnOut183= MEMEnIn1[83:83];
assign MEMRWEnOut183= MEMRWEnIn1[83:83];
assign MEMDataOut83= mLocalDataIn[2687:2656];
assign mLocalDataOut[2687:2656] = MEMDataIn83;
assign MEMAddrOut183= MEMAddrIn1[503:498];
assign MEMEnOut184= MEMEnIn1[84:84];
assign MEMRWEnOut184= MEMRWEnIn1[84:84];
assign MEMDataOut84= mLocalDataIn[2719:2688];
assign mLocalDataOut[2719:2688] = MEMDataIn84;
assign MEMAddrOut184= MEMAddrIn1[509:504];
assign MEMEnOut185= MEMEnIn1[85:85];
assign MEMRWEnOut185= MEMRWEnIn1[85:85];
assign MEMDataOut85= mLocalDataIn[2751:2720];
assign mLocalDataOut[2751:2720] = MEMDataIn85;
assign MEMAddrOut185= MEMAddrIn1[515:510];
assign MEMEnOut186= MEMEnIn1[86:86];
assign MEMRWEnOut186= MEMRWEnIn1[86:86];
assign MEMDataOut86= mLocalDataIn[2783:2752];
assign mLocalDataOut[2783:2752] = MEMDataIn86;
assign MEMAddrOut186= MEMAddrIn1[521:516];
assign MEMEnOut187= MEMEnIn1[87:87];
assign MEMRWEnOut187= MEMRWEnIn1[87:87];
assign MEMDataOut87= mLocalDataIn[2815:2784];
assign mLocalDataOut[2815:2784] = MEMDataIn87;
assign MEMAddrOut187= MEMAddrIn1[527:522];
assign MEMEnOut188= MEMEnIn1[88:88];
assign MEMRWEnOut188= MEMRWEnIn1[88:88];
assign MEMDataOut88= mLocalDataIn[2847:2816];
assign mLocalDataOut[2847:2816] = MEMDataIn88;
assign MEMAddrOut188= MEMAddrIn1[533:528];
assign MEMEnOut189= MEMEnIn1[89:89];
assign MEMRWEnOut189= MEMRWEnIn1[89:89];
assign MEMDataOut89= mLocalDataIn[2879:2848];
assign mLocalDataOut[2879:2848] = MEMDataIn89;
assign MEMAddrOut189= MEMAddrIn1[539:534];
assign MEMEnOut190= MEMEnIn1[90:90];
assign MEMRWEnOut190= MEMRWEnIn1[90:90];
assign MEMDataOut90= mLocalDataIn[2911:2880];
assign mLocalDataOut[2911:2880] = MEMDataIn90;
assign MEMAddrOut190= MEMAddrIn1[545:540];
assign MEMEnOut191= MEMEnIn1[91:91];
assign MEMRWEnOut191= MEMRWEnIn1[91:91];
assign MEMDataOut91= mLocalDataIn[2943:2912];
assign mLocalDataOut[2943:2912] = MEMDataIn91;
assign MEMAddrOut191= MEMAddrIn1[551:546];
assign MEMEnOut192= MEMEnIn1[92:92];
assign MEMRWEnOut192= MEMRWEnIn1[92:92];
assign MEMDataOut92= mLocalDataIn[2975:2944];
assign mLocalDataOut[2975:2944] = MEMDataIn92;
assign MEMAddrOut192= MEMAddrIn1[557:552];
assign MEMEnOut193= MEMEnIn1[93:93];
assign MEMRWEnOut193= MEMRWEnIn1[93:93];
assign MEMDataOut93= mLocalDataIn[3007:2976];
assign mLocalDataOut[3007:2976] = MEMDataIn93;
assign MEMAddrOut193= MEMAddrIn1[563:558];
assign MEMEnOut194= MEMEnIn1[94:94];
assign MEMRWEnOut194= MEMRWEnIn1[94:94];
assign MEMDataOut94= mLocalDataIn[3039:3008];
assign mLocalDataOut[3039:3008] = MEMDataIn94;
assign MEMAddrOut194= MEMAddrIn1[569:564];
assign MEMEnOut195= MEMEnIn1[95:95];
assign MEMRWEnOut195= MEMRWEnIn1[95:95];
assign MEMDataOut95= mLocalDataIn[3071:3040];
assign mLocalDataOut[3071:3040] = MEMDataIn95;
assign MEMAddrOut195= MEMAddrIn1[575:570];
assign MEMEnOut196= MEMEnIn1[96:96];
assign MEMRWEnOut196= MEMRWEnIn1[96:96];
assign MEMDataOut96= mLocalDataIn[3103:3072];
assign mLocalDataOut[3103:3072] = MEMDataIn96;
assign MEMAddrOut196= MEMAddrIn1[581:576];
assign MEMEnOut197= MEMEnIn1[97:97];
assign MEMRWEnOut197= MEMRWEnIn1[97:97];
assign MEMDataOut97= mLocalDataIn[3135:3104];
assign mLocalDataOut[3135:3104] = MEMDataIn97;
assign MEMAddrOut197= MEMAddrIn1[587:582];
assign MEMEnOut198= MEMEnIn1[98:98];
assign MEMRWEnOut198= MEMRWEnIn1[98:98];
assign MEMDataOut98= mLocalDataIn[3167:3136];
assign mLocalDataOut[3167:3136] = MEMDataIn98;
assign MEMAddrOut198= MEMAddrIn1[593:588];
assign MEMEnOut199= MEMEnIn1[99:99];
assign MEMRWEnOut199= MEMRWEnIn1[99:99];
assign MEMDataOut99= mLocalDataIn[3199:3168];
assign mLocalDataOut[3199:3168] = MEMDataIn99;
assign MEMAddrOut199= MEMAddrIn1[599:594];
assign MEMEnOut1100= MEMEnIn1[100:100];
assign MEMRWEnOut1100= MEMRWEnIn1[100:100];
assign MEMDataOut100= mLocalDataIn[3231:3200];
assign mLocalDataOut[3231:3200] = MEMDataIn100;
assign MEMAddrOut1100= MEMAddrIn1[605:600];
assign MEMEnOut1101= MEMEnIn1[101:101];
assign MEMRWEnOut1101= MEMRWEnIn1[101:101];
assign MEMDataOut101= mLocalDataIn[3263:3232];
assign mLocalDataOut[3263:3232] = MEMDataIn101;
assign MEMAddrOut1101= MEMAddrIn1[611:606];
assign MEMEnOut1102= MEMEnIn1[102:102];
assign MEMRWEnOut1102= MEMRWEnIn1[102:102];
assign MEMDataOut102= mLocalDataIn[3295:3264];
assign mLocalDataOut[3295:3264] = MEMDataIn102;
assign MEMAddrOut1102= MEMAddrIn1[617:612];
assign MEMEnOut1103= MEMEnIn1[103:103];
assign MEMRWEnOut1103= MEMRWEnIn1[103:103];
assign MEMDataOut103= mLocalDataIn[3327:3296];
assign mLocalDataOut[3327:3296] = MEMDataIn103;
assign MEMAddrOut1103= MEMAddrIn1[623:618];
assign MEMEnOut1104= MEMEnIn1[104:104];
assign MEMRWEnOut1104= MEMRWEnIn1[104:104];
assign MEMDataOut104= mLocalDataIn[3359:3328];
assign mLocalDataOut[3359:3328] = MEMDataIn104;
assign MEMAddrOut1104= MEMAddrIn1[629:624];
assign MEMEnOut1105= MEMEnIn1[105:105];
assign MEMRWEnOut1105= MEMRWEnIn1[105:105];
assign MEMDataOut105= mLocalDataIn[3391:3360];
assign mLocalDataOut[3391:3360] = MEMDataIn105;
assign MEMAddrOut1105= MEMAddrIn1[635:630];
assign MEMEnOut1106= MEMEnIn1[106:106];
assign MEMRWEnOut1106= MEMRWEnIn1[106:106];
assign MEMDataOut106= mLocalDataIn[3423:3392];
assign mLocalDataOut[3423:3392] = MEMDataIn106;
assign MEMAddrOut1106= MEMAddrIn1[641:636];
assign MEMEnOut1107= MEMEnIn1[107:107];
assign MEMRWEnOut1107= MEMRWEnIn1[107:107];
assign MEMDataOut107= mLocalDataIn[3455:3424];
assign mLocalDataOut[3455:3424] = MEMDataIn107;
assign MEMAddrOut1107= MEMAddrIn1[647:642];
output [38:0] IMEMDataOut;
input [38:0] IMEMDataIn;
assign IMEMDataOut = mILocalDataIn;
assign mILocalDataOut = IMEMDataIn;
assign IMEMEnOut1 = IMEMEnIn1;
assign IMEMRWEnOut1 = IMEMRWEnIn1;
assign IMEMAddrOut1 = IMEMAddrIn1;
output MEMEnOut20;
output MEMRWEnOut20;
output [5:0] MEMAddrOut20;
output MEMEnOut21;
output MEMRWEnOut21;
output [5:0] MEMAddrOut21;
output MEMEnOut22;
output MEMRWEnOut22;
output [5:0] MEMAddrOut22;
output MEMEnOut23;
output MEMRWEnOut23;
output [5:0] MEMAddrOut23;
output MEMEnOut24;
output MEMRWEnOut24;
output [5:0] MEMAddrOut24;
output MEMEnOut25;
output MEMRWEnOut25;
output [5:0] MEMAddrOut25;
output MEMEnOut26;
output MEMRWEnOut26;
output [5:0] MEMAddrOut26;
output MEMEnOut27;
output MEMRWEnOut27;
output [5:0] MEMAddrOut27;
output MEMEnOut28;
output MEMRWEnOut28;
output [5:0] MEMAddrOut28;
output MEMEnOut29;
output MEMRWEnOut29;
output [5:0] MEMAddrOut29;
output MEMEnOut210;
output MEMRWEnOut210;
output [5:0] MEMAddrOut210;
output MEMEnOut211;
output MEMRWEnOut211;
output [5:0] MEMAddrOut211;
output MEMEnOut212;
output MEMRWEnOut212;
output [5:0] MEMAddrOut212;
output MEMEnOut213;
output MEMRWEnOut213;
output [5:0] MEMAddrOut213;
output MEMEnOut214;
output MEMRWEnOut214;
output [5:0] MEMAddrOut214;
output MEMEnOut215;
output MEMRWEnOut215;
output [5:0] MEMAddrOut215;
output MEMEnOut216;
output MEMRWEnOut216;
output [5:0] MEMAddrOut216;
output MEMEnOut217;
output MEMRWEnOut217;
output [5:0] MEMAddrOut217;
output MEMEnOut218;
output MEMRWEnOut218;
output [5:0] MEMAddrOut218;
output MEMEnOut219;
output MEMRWEnOut219;
output [5:0] MEMAddrOut219;
output MEMEnOut220;
output MEMRWEnOut220;
output [5:0] MEMAddrOut220;
output MEMEnOut221;
output MEMRWEnOut221;
output [5:0] MEMAddrOut221;
output MEMEnOut222;
output MEMRWEnOut222;
output [5:0] MEMAddrOut222;
output MEMEnOut223;
output MEMRWEnOut223;
output [5:0] MEMAddrOut223;
output MEMEnOut224;
output MEMRWEnOut224;
output [5:0] MEMAddrOut224;
output MEMEnOut225;
output MEMRWEnOut225;
output [5:0] MEMAddrOut225;
output MEMEnOut226;
output MEMRWEnOut226;
output [5:0] MEMAddrOut226;
output MEMEnOut227;
output MEMRWEnOut227;
output [5:0] MEMAddrOut227;
output MEMEnOut228;
output MEMRWEnOut228;
output [5:0] MEMAddrOut228;
output MEMEnOut229;
output MEMRWEnOut229;
output [5:0] MEMAddrOut229;
output MEMEnOut230;
output MEMRWEnOut230;
output [5:0] MEMAddrOut230;
output MEMEnOut231;
output MEMRWEnOut231;
output [5:0] MEMAddrOut231;
output MEMEnOut232;
output MEMRWEnOut232;
output [5:0] MEMAddrOut232;
output MEMEnOut233;
output MEMRWEnOut233;
output [5:0] MEMAddrOut233;
output MEMEnOut234;
output MEMRWEnOut234;
output [5:0] MEMAddrOut234;
output MEMEnOut235;
output MEMRWEnOut235;
output [5:0] MEMAddrOut235;
output MEMEnOut236;
output MEMRWEnOut236;
output [5:0] MEMAddrOut236;
output MEMEnOut237;
output MEMRWEnOut237;
output [5:0] MEMAddrOut237;
output MEMEnOut238;
output MEMRWEnOut238;
output [5:0] MEMAddrOut238;
output MEMEnOut239;
output MEMRWEnOut239;
output [5:0] MEMAddrOut239;
output MEMEnOut240;
output MEMRWEnOut240;
output [5:0] MEMAddrOut240;
output MEMEnOut241;
output MEMRWEnOut241;
output [5:0] MEMAddrOut241;
output MEMEnOut242;
output MEMRWEnOut242;
output [5:0] MEMAddrOut242;
output MEMEnOut243;
output MEMRWEnOut243;
output [5:0] MEMAddrOut243;
output MEMEnOut244;
output MEMRWEnOut244;
output [5:0] MEMAddrOut244;
output MEMEnOut245;
output MEMRWEnOut245;
output [5:0] MEMAddrOut245;
output MEMEnOut246;
output MEMRWEnOut246;
output [5:0] MEMAddrOut246;
output MEMEnOut247;
output MEMRWEnOut247;
output [5:0] MEMAddrOut247;
output MEMEnOut248;
output MEMRWEnOut248;
output [5:0] MEMAddrOut248;
output MEMEnOut249;
output MEMRWEnOut249;
output [5:0] MEMAddrOut249;
output MEMEnOut250;
output MEMRWEnOut250;
output [5:0] MEMAddrOut250;
output MEMEnOut251;
output MEMRWEnOut251;
output [5:0] MEMAddrOut251;
output MEMEnOut252;
output MEMRWEnOut252;
output [5:0] MEMAddrOut252;
output MEMEnOut253;
output MEMRWEnOut253;
output [5:0] MEMAddrOut253;
output MEMEnOut254;
output MEMRWEnOut254;
output [5:0] MEMAddrOut254;
output MEMEnOut255;
output MEMRWEnOut255;
output [5:0] MEMAddrOut255;
output MEMEnOut256;
output MEMRWEnOut256;
output [5:0] MEMAddrOut256;
output MEMEnOut257;
output MEMRWEnOut257;
output [5:0] MEMAddrOut257;
output MEMEnOut258;
output MEMRWEnOut258;
output [5:0] MEMAddrOut258;
output MEMEnOut259;
output MEMRWEnOut259;
output [5:0] MEMAddrOut259;
output MEMEnOut260;
output MEMRWEnOut260;
output [5:0] MEMAddrOut260;
output MEMEnOut261;
output MEMRWEnOut261;
output [5:0] MEMAddrOut261;
output MEMEnOut262;
output MEMRWEnOut262;
output [5:0] MEMAddrOut262;
output MEMEnOut263;
output MEMRWEnOut263;
output [5:0] MEMAddrOut263;
output MEMEnOut264;
output MEMRWEnOut264;
output [5:0] MEMAddrOut264;
output MEMEnOut265;
output MEMRWEnOut265;
output [5:0] MEMAddrOut265;
output MEMEnOut266;
output MEMRWEnOut266;
output [5:0] MEMAddrOut266;
output MEMEnOut267;
output MEMRWEnOut267;
output [5:0] MEMAddrOut267;
output MEMEnOut268;
output MEMRWEnOut268;
output [5:0] MEMAddrOut268;
output MEMEnOut269;
output MEMRWEnOut269;
output [5:0] MEMAddrOut269;
output MEMEnOut270;
output MEMRWEnOut270;
output [5:0] MEMAddrOut270;
output MEMEnOut271;
output MEMRWEnOut271;
output [5:0] MEMAddrOut271;
output MEMEnOut272;
output MEMRWEnOut272;
output [5:0] MEMAddrOut272;
output MEMEnOut273;
output MEMRWEnOut273;
output [5:0] MEMAddrOut273;
output MEMEnOut274;
output MEMRWEnOut274;
output [5:0] MEMAddrOut274;
output MEMEnOut275;
output MEMRWEnOut275;
output [5:0] MEMAddrOut275;
output MEMEnOut276;
output MEMRWEnOut276;
output [5:0] MEMAddrOut276;
output MEMEnOut277;
output MEMRWEnOut277;
output [5:0] MEMAddrOut277;
output MEMEnOut278;
output MEMRWEnOut278;
output [5:0] MEMAddrOut278;
output MEMEnOut279;
output MEMRWEnOut279;
output [5:0] MEMAddrOut279;
output MEMEnOut280;
output MEMRWEnOut280;
output [5:0] MEMAddrOut280;
output MEMEnOut281;
output MEMRWEnOut281;
output [5:0] MEMAddrOut281;
output MEMEnOut282;
output MEMRWEnOut282;
output [5:0] MEMAddrOut282;
output MEMEnOut283;
output MEMRWEnOut283;
output [5:0] MEMAddrOut283;
output MEMEnOut284;
output MEMRWEnOut284;
output [5:0] MEMAddrOut284;
output MEMEnOut285;
output MEMRWEnOut285;
output [5:0] MEMAddrOut285;
output MEMEnOut286;
output MEMRWEnOut286;
output [5:0] MEMAddrOut286;
output MEMEnOut287;
output MEMRWEnOut287;
output [5:0] MEMAddrOut287;
output MEMEnOut288;
output MEMRWEnOut288;
output [5:0] MEMAddrOut288;
output MEMEnOut289;
output MEMRWEnOut289;
output [5:0] MEMAddrOut289;
output MEMEnOut290;
output MEMRWEnOut290;
output [5:0] MEMAddrOut290;
output MEMEnOut291;
output MEMRWEnOut291;
output [5:0] MEMAddrOut291;
output MEMEnOut292;
output MEMRWEnOut292;
output [5:0] MEMAddrOut292;
output MEMEnOut293;
output MEMRWEnOut293;
output [5:0] MEMAddrOut293;
output MEMEnOut294;
output MEMRWEnOut294;
output [5:0] MEMAddrOut294;
output MEMEnOut295;
output MEMRWEnOut295;
output [5:0] MEMAddrOut295;
output MEMEnOut296;
output MEMRWEnOut296;
output [5:0] MEMAddrOut296;
output MEMEnOut297;
output MEMRWEnOut297;
output [5:0] MEMAddrOut297;
output MEMEnOut298;
output MEMRWEnOut298;
output [5:0] MEMAddrOut298;
output MEMEnOut299;
output MEMRWEnOut299;
output [5:0] MEMAddrOut299;
output MEMEnOut2100;
output MEMRWEnOut2100;
output [5:0] MEMAddrOut2100;
output MEMEnOut2101;
output MEMRWEnOut2101;
output [5:0] MEMAddrOut2101;
output MEMEnOut2102;
output MEMRWEnOut2102;
output [5:0] MEMAddrOut2102;
output MEMEnOut2103;
output MEMRWEnOut2103;
output [5:0] MEMAddrOut2103;
output MEMEnOut2104;
output MEMRWEnOut2104;
output [5:0] MEMAddrOut2104;
output MEMEnOut2105;
output MEMRWEnOut2105;
output [5:0] MEMAddrOut2105;
output MEMEnOut2106;
output MEMRWEnOut2106;
output [5:0] MEMAddrOut2106;
output MEMEnOut2107;
output MEMRWEnOut2107;
output [5:0] MEMAddrOut2107;
assign MEMEnOut20= MEMEnIn2[0:0];
assign MEMRWEnOut20= MEMRWEnIn2[0:0];
assign MEMAddrOut20= MEMAddrIn2[5:0];
assign MEMEnOut21= MEMEnIn2[1:1];
assign MEMRWEnOut21= MEMRWEnIn2[1:1];
assign MEMAddrOut21= MEMAddrIn2[11:6];
assign MEMEnOut22= MEMEnIn2[2:2];
assign MEMRWEnOut22= MEMRWEnIn2[2:2];
assign MEMAddrOut22= MEMAddrIn2[17:12];
assign MEMEnOut23= MEMEnIn2[3:3];
assign MEMRWEnOut23= MEMRWEnIn2[3:3];
assign MEMAddrOut23= MEMAddrIn2[23:18];
assign MEMEnOut24= MEMEnIn2[4:4];
assign MEMRWEnOut24= MEMRWEnIn2[4:4];
assign MEMAddrOut24= MEMAddrIn2[29:24];
assign MEMEnOut25= MEMEnIn2[5:5];
assign MEMRWEnOut25= MEMRWEnIn2[5:5];
assign MEMAddrOut25= MEMAddrIn2[35:30];
assign MEMEnOut26= MEMEnIn2[6:6];
assign MEMRWEnOut26= MEMRWEnIn2[6:6];
assign MEMAddrOut26= MEMAddrIn2[41:36];
assign MEMEnOut27= MEMEnIn2[7:7];
assign MEMRWEnOut27= MEMRWEnIn2[7:7];
assign MEMAddrOut27= MEMAddrIn2[47:42];
assign MEMEnOut28= MEMEnIn2[8:8];
assign MEMRWEnOut28= MEMRWEnIn2[8:8];
assign MEMAddrOut28= MEMAddrIn2[53:48];
assign MEMEnOut29= MEMEnIn2[9:9];
assign MEMRWEnOut29= MEMRWEnIn2[9:9];
assign MEMAddrOut29= MEMAddrIn2[59:54];
assign MEMEnOut210= MEMEnIn2[10:10];
assign MEMRWEnOut210= MEMRWEnIn2[10:10];
assign MEMAddrOut210= MEMAddrIn2[65:60];
assign MEMEnOut211= MEMEnIn2[11:11];
assign MEMRWEnOut211= MEMRWEnIn2[11:11];
assign MEMAddrOut211= MEMAddrIn2[71:66];
assign MEMEnOut212= MEMEnIn2[12:12];
assign MEMRWEnOut212= MEMRWEnIn2[12:12];
assign MEMAddrOut212= MEMAddrIn2[77:72];
assign MEMEnOut213= MEMEnIn2[13:13];
assign MEMRWEnOut213= MEMRWEnIn2[13:13];
assign MEMAddrOut213= MEMAddrIn2[83:78];
assign MEMEnOut214= MEMEnIn2[14:14];
assign MEMRWEnOut214= MEMRWEnIn2[14:14];
assign MEMAddrOut214= MEMAddrIn2[89:84];
assign MEMEnOut215= MEMEnIn2[15:15];
assign MEMRWEnOut215= MEMRWEnIn2[15:15];
assign MEMAddrOut215= MEMAddrIn2[95:90];
assign MEMEnOut216= MEMEnIn2[16:16];
assign MEMRWEnOut216= MEMRWEnIn2[16:16];
assign MEMAddrOut216= MEMAddrIn2[101:96];
assign MEMEnOut217= MEMEnIn2[17:17];
assign MEMRWEnOut217= MEMRWEnIn2[17:17];
assign MEMAddrOut217= MEMAddrIn2[107:102];
assign MEMEnOut218= MEMEnIn2[18:18];
assign MEMRWEnOut218= MEMRWEnIn2[18:18];
assign MEMAddrOut218= MEMAddrIn2[113:108];
assign MEMEnOut219= MEMEnIn2[19:19];
assign MEMRWEnOut219= MEMRWEnIn2[19:19];
assign MEMAddrOut219= MEMAddrIn2[119:114];
assign MEMEnOut220= MEMEnIn2[20:20];
assign MEMRWEnOut220= MEMRWEnIn2[20:20];
assign MEMAddrOut220= MEMAddrIn2[125:120];
assign MEMEnOut221= MEMEnIn2[21:21];
assign MEMRWEnOut221= MEMRWEnIn2[21:21];
assign MEMAddrOut221= MEMAddrIn2[131:126];
assign MEMEnOut222= MEMEnIn2[22:22];
assign MEMRWEnOut222= MEMRWEnIn2[22:22];
assign MEMAddrOut222= MEMAddrIn2[137:132];
assign MEMEnOut223= MEMEnIn2[23:23];
assign MEMRWEnOut223= MEMRWEnIn2[23:23];
assign MEMAddrOut223= MEMAddrIn2[143:138];
assign MEMEnOut224= MEMEnIn2[24:24];
assign MEMRWEnOut224= MEMRWEnIn2[24:24];
assign MEMAddrOut224= MEMAddrIn2[149:144];
assign MEMEnOut225= MEMEnIn2[25:25];
assign MEMRWEnOut225= MEMRWEnIn2[25:25];
assign MEMAddrOut225= MEMAddrIn2[155:150];
assign MEMEnOut226= MEMEnIn2[26:26];
assign MEMRWEnOut226= MEMRWEnIn2[26:26];
assign MEMAddrOut226= MEMAddrIn2[161:156];
assign MEMEnOut227= MEMEnIn2[27:27];
assign MEMRWEnOut227= MEMRWEnIn2[27:27];
assign MEMAddrOut227= MEMAddrIn2[167:162];
assign MEMEnOut228= MEMEnIn2[28:28];
assign MEMRWEnOut228= MEMRWEnIn2[28:28];
assign MEMAddrOut228= MEMAddrIn2[173:168];
assign MEMEnOut229= MEMEnIn2[29:29];
assign MEMRWEnOut229= MEMRWEnIn2[29:29];
assign MEMAddrOut229= MEMAddrIn2[179:174];
assign MEMEnOut230= MEMEnIn2[30:30];
assign MEMRWEnOut230= MEMRWEnIn2[30:30];
assign MEMAddrOut230= MEMAddrIn2[185:180];
assign MEMEnOut231= MEMEnIn2[31:31];
assign MEMRWEnOut231= MEMRWEnIn2[31:31];
assign MEMAddrOut231= MEMAddrIn2[191:186];
assign MEMEnOut232= MEMEnIn2[32:32];
assign MEMRWEnOut232= MEMRWEnIn2[32:32];
assign MEMAddrOut232= MEMAddrIn2[197:192];
assign MEMEnOut233= MEMEnIn2[33:33];
assign MEMRWEnOut233= MEMRWEnIn2[33:33];
assign MEMAddrOut233= MEMAddrIn2[203:198];
assign MEMEnOut234= MEMEnIn2[34:34];
assign MEMRWEnOut234= MEMRWEnIn2[34:34];
assign MEMAddrOut234= MEMAddrIn2[209:204];
assign MEMEnOut235= MEMEnIn2[35:35];
assign MEMRWEnOut235= MEMRWEnIn2[35:35];
assign MEMAddrOut235= MEMAddrIn2[215:210];
assign MEMEnOut236= MEMEnIn2[36:36];
assign MEMRWEnOut236= MEMRWEnIn2[36:36];
assign MEMAddrOut236= MEMAddrIn2[221:216];
assign MEMEnOut237= MEMEnIn2[37:37];
assign MEMRWEnOut237= MEMRWEnIn2[37:37];
assign MEMAddrOut237= MEMAddrIn2[227:222];
assign MEMEnOut238= MEMEnIn2[38:38];
assign MEMRWEnOut238= MEMRWEnIn2[38:38];
assign MEMAddrOut238= MEMAddrIn2[233:228];
assign MEMEnOut239= MEMEnIn2[39:39];
assign MEMRWEnOut239= MEMRWEnIn2[39:39];
assign MEMAddrOut239= MEMAddrIn2[239:234];
assign MEMEnOut240= MEMEnIn2[40:40];
assign MEMRWEnOut240= MEMRWEnIn2[40:40];
assign MEMAddrOut240= MEMAddrIn2[245:240];
assign MEMEnOut241= MEMEnIn2[41:41];
assign MEMRWEnOut241= MEMRWEnIn2[41:41];
assign MEMAddrOut241= MEMAddrIn2[251:246];
assign MEMEnOut242= MEMEnIn2[42:42];
assign MEMRWEnOut242= MEMRWEnIn2[42:42];
assign MEMAddrOut242= MEMAddrIn2[257:252];
assign MEMEnOut243= MEMEnIn2[43:43];
assign MEMRWEnOut243= MEMRWEnIn2[43:43];
assign MEMAddrOut243= MEMAddrIn2[263:258];
assign MEMEnOut244= MEMEnIn2[44:44];
assign MEMRWEnOut244= MEMRWEnIn2[44:44];
assign MEMAddrOut244= MEMAddrIn2[269:264];
assign MEMEnOut245= MEMEnIn2[45:45];
assign MEMRWEnOut245= MEMRWEnIn2[45:45];
assign MEMAddrOut245= MEMAddrIn2[275:270];
assign MEMEnOut246= MEMEnIn2[46:46];
assign MEMRWEnOut246= MEMRWEnIn2[46:46];
assign MEMAddrOut246= MEMAddrIn2[281:276];
assign MEMEnOut247= MEMEnIn2[47:47];
assign MEMRWEnOut247= MEMRWEnIn2[47:47];
assign MEMAddrOut247= MEMAddrIn2[287:282];
assign MEMEnOut248= MEMEnIn2[48:48];
assign MEMRWEnOut248= MEMRWEnIn2[48:48];
assign MEMAddrOut248= MEMAddrIn2[293:288];
assign MEMEnOut249= MEMEnIn2[49:49];
assign MEMRWEnOut249= MEMRWEnIn2[49:49];
assign MEMAddrOut249= MEMAddrIn2[299:294];
assign MEMEnOut250= MEMEnIn2[50:50];
assign MEMRWEnOut250= MEMRWEnIn2[50:50];
assign MEMAddrOut250= MEMAddrIn2[305:300];
assign MEMEnOut251= MEMEnIn2[51:51];
assign MEMRWEnOut251= MEMRWEnIn2[51:51];
assign MEMAddrOut251= MEMAddrIn2[311:306];
assign MEMEnOut252= MEMEnIn2[52:52];
assign MEMRWEnOut252= MEMRWEnIn2[52:52];
assign MEMAddrOut252= MEMAddrIn2[317:312];
assign MEMEnOut253= MEMEnIn2[53:53];
assign MEMRWEnOut253= MEMRWEnIn2[53:53];
assign MEMAddrOut253= MEMAddrIn2[323:318];
assign MEMEnOut254= MEMEnIn2[54:54];
assign MEMRWEnOut254= MEMRWEnIn2[54:54];
assign MEMAddrOut254= MEMAddrIn2[329:324];
assign MEMEnOut255= MEMEnIn2[55:55];
assign MEMRWEnOut255= MEMRWEnIn2[55:55];
assign MEMAddrOut255= MEMAddrIn2[335:330];
assign MEMEnOut256= MEMEnIn2[56:56];
assign MEMRWEnOut256= MEMRWEnIn2[56:56];
assign MEMAddrOut256= MEMAddrIn2[341:336];
assign MEMEnOut257= MEMEnIn2[57:57];
assign MEMRWEnOut257= MEMRWEnIn2[57:57];
assign MEMAddrOut257= MEMAddrIn2[347:342];
assign MEMEnOut258= MEMEnIn2[58:58];
assign MEMRWEnOut258= MEMRWEnIn2[58:58];
assign MEMAddrOut258= MEMAddrIn2[353:348];
assign MEMEnOut259= MEMEnIn2[59:59];
assign MEMRWEnOut259= MEMRWEnIn2[59:59];
assign MEMAddrOut259= MEMAddrIn2[359:354];
assign MEMEnOut260= MEMEnIn2[60:60];
assign MEMRWEnOut260= MEMRWEnIn2[60:60];
assign MEMAddrOut260= MEMAddrIn2[365:360];
assign MEMEnOut261= MEMEnIn2[61:61];
assign MEMRWEnOut261= MEMRWEnIn2[61:61];
assign MEMAddrOut261= MEMAddrIn2[371:366];
assign MEMEnOut262= MEMEnIn2[62:62];
assign MEMRWEnOut262= MEMRWEnIn2[62:62];
assign MEMAddrOut262= MEMAddrIn2[377:372];
assign MEMEnOut263= MEMEnIn2[63:63];
assign MEMRWEnOut263= MEMRWEnIn2[63:63];
assign MEMAddrOut263= MEMAddrIn2[383:378];
assign MEMEnOut264= MEMEnIn2[64:64];
assign MEMRWEnOut264= MEMRWEnIn2[64:64];
assign MEMAddrOut264= MEMAddrIn2[389:384];
assign MEMEnOut265= MEMEnIn2[65:65];
assign MEMRWEnOut265= MEMRWEnIn2[65:65];
assign MEMAddrOut265= MEMAddrIn2[395:390];
assign MEMEnOut266= MEMEnIn2[66:66];
assign MEMRWEnOut266= MEMRWEnIn2[66:66];
assign MEMAddrOut266= MEMAddrIn2[401:396];
assign MEMEnOut267= MEMEnIn2[67:67];
assign MEMRWEnOut267= MEMRWEnIn2[67:67];
assign MEMAddrOut267= MEMAddrIn2[407:402];
assign MEMEnOut268= MEMEnIn2[68:68];
assign MEMRWEnOut268= MEMRWEnIn2[68:68];
assign MEMAddrOut268= MEMAddrIn2[413:408];
assign MEMEnOut269= MEMEnIn2[69:69];
assign MEMRWEnOut269= MEMRWEnIn2[69:69];
assign MEMAddrOut269= MEMAddrIn2[419:414];
assign MEMEnOut270= MEMEnIn2[70:70];
assign MEMRWEnOut270= MEMRWEnIn2[70:70];
assign MEMAddrOut270= MEMAddrIn2[425:420];
assign MEMEnOut271= MEMEnIn2[71:71];
assign MEMRWEnOut271= MEMRWEnIn2[71:71];
assign MEMAddrOut271= MEMAddrIn2[431:426];
assign MEMEnOut272= MEMEnIn2[72:72];
assign MEMRWEnOut272= MEMRWEnIn2[72:72];
assign MEMAddrOut272= MEMAddrIn2[437:432];
assign MEMEnOut273= MEMEnIn2[73:73];
assign MEMRWEnOut273= MEMRWEnIn2[73:73];
assign MEMAddrOut273= MEMAddrIn2[443:438];
assign MEMEnOut274= MEMEnIn2[74:74];
assign MEMRWEnOut274= MEMRWEnIn2[74:74];
assign MEMAddrOut274= MEMAddrIn2[449:444];
assign MEMEnOut275= MEMEnIn2[75:75];
assign MEMRWEnOut275= MEMRWEnIn2[75:75];
assign MEMAddrOut275= MEMAddrIn2[455:450];
assign MEMEnOut276= MEMEnIn2[76:76];
assign MEMRWEnOut276= MEMRWEnIn2[76:76];
assign MEMAddrOut276= MEMAddrIn2[461:456];
assign MEMEnOut277= MEMEnIn2[77:77];
assign MEMRWEnOut277= MEMRWEnIn2[77:77];
assign MEMAddrOut277= MEMAddrIn2[467:462];
assign MEMEnOut278= MEMEnIn2[78:78];
assign MEMRWEnOut278= MEMRWEnIn2[78:78];
assign MEMAddrOut278= MEMAddrIn2[473:468];
assign MEMEnOut279= MEMEnIn2[79:79];
assign MEMRWEnOut279= MEMRWEnIn2[79:79];
assign MEMAddrOut279= MEMAddrIn2[479:474];
assign MEMEnOut280= MEMEnIn2[80:80];
assign MEMRWEnOut280= MEMRWEnIn2[80:80];
assign MEMAddrOut280= MEMAddrIn2[485:480];
assign MEMEnOut281= MEMEnIn2[81:81];
assign MEMRWEnOut281= MEMRWEnIn2[81:81];
assign MEMAddrOut281= MEMAddrIn2[491:486];
assign MEMEnOut282= MEMEnIn2[82:82];
assign MEMRWEnOut282= MEMRWEnIn2[82:82];
assign MEMAddrOut282= MEMAddrIn2[497:492];
assign MEMEnOut283= MEMEnIn2[83:83];
assign MEMRWEnOut283= MEMRWEnIn2[83:83];
assign MEMAddrOut283= MEMAddrIn2[503:498];
assign MEMEnOut284= MEMEnIn2[84:84];
assign MEMRWEnOut284= MEMRWEnIn2[84:84];
assign MEMAddrOut284= MEMAddrIn2[509:504];
assign MEMEnOut285= MEMEnIn2[85:85];
assign MEMRWEnOut285= MEMRWEnIn2[85:85];
assign MEMAddrOut285= MEMAddrIn2[515:510];
assign MEMEnOut286= MEMEnIn2[86:86];
assign MEMRWEnOut286= MEMRWEnIn2[86:86];
assign MEMAddrOut286= MEMAddrIn2[521:516];
assign MEMEnOut287= MEMEnIn2[87:87];
assign MEMRWEnOut287= MEMRWEnIn2[87:87];
assign MEMAddrOut287= MEMAddrIn2[527:522];
assign MEMEnOut288= MEMEnIn2[88:88];
assign MEMRWEnOut288= MEMRWEnIn2[88:88];
assign MEMAddrOut288= MEMAddrIn2[533:528];
assign MEMEnOut289= MEMEnIn2[89:89];
assign MEMRWEnOut289= MEMRWEnIn2[89:89];
assign MEMAddrOut289= MEMAddrIn2[539:534];
assign MEMEnOut290= MEMEnIn2[90:90];
assign MEMRWEnOut290= MEMRWEnIn2[90:90];
assign MEMAddrOut290= MEMAddrIn2[545:540];
assign MEMEnOut291= MEMEnIn2[91:91];
assign MEMRWEnOut291= MEMRWEnIn2[91:91];
assign MEMAddrOut291= MEMAddrIn2[551:546];
assign MEMEnOut292= MEMEnIn2[92:92];
assign MEMRWEnOut292= MEMRWEnIn2[92:92];
assign MEMAddrOut292= MEMAddrIn2[557:552];
assign MEMEnOut293= MEMEnIn2[93:93];
assign MEMRWEnOut293= MEMRWEnIn2[93:93];
assign MEMAddrOut293= MEMAddrIn2[563:558];
assign MEMEnOut294= MEMEnIn2[94:94];
assign MEMRWEnOut294= MEMRWEnIn2[94:94];
assign MEMAddrOut294= MEMAddrIn2[569:564];
assign MEMEnOut295= MEMEnIn2[95:95];
assign MEMRWEnOut295= MEMRWEnIn2[95:95];
assign MEMAddrOut295= MEMAddrIn2[575:570];
assign MEMEnOut296= MEMEnIn2[96:96];
assign MEMRWEnOut296= MEMRWEnIn2[96:96];
assign MEMAddrOut296= MEMAddrIn2[581:576];
assign MEMEnOut297= MEMEnIn2[97:97];
assign MEMRWEnOut297= MEMRWEnIn2[97:97];
assign MEMAddrOut297= MEMAddrIn2[587:582];
assign MEMEnOut298= MEMEnIn2[98:98];
assign MEMRWEnOut298= MEMRWEnIn2[98:98];
assign MEMAddrOut298= MEMAddrIn2[593:588];
assign MEMEnOut299= MEMEnIn2[99:99];
assign MEMRWEnOut299= MEMRWEnIn2[99:99];
assign MEMAddrOut299= MEMAddrIn2[599:594];
assign MEMEnOut2100= MEMEnIn2[100:100];
assign MEMRWEnOut2100= MEMRWEnIn2[100:100];
assign MEMAddrOut2100= MEMAddrIn2[605:600];
assign MEMEnOut2101= MEMEnIn2[101:101];
assign MEMRWEnOut2101= MEMRWEnIn2[101:101];
assign MEMAddrOut2101= MEMAddrIn2[611:606];
assign MEMEnOut2102= MEMEnIn2[102:102];
assign MEMRWEnOut2102= MEMRWEnIn2[102:102];
assign MEMAddrOut2102= MEMAddrIn2[617:612];
assign MEMEnOut2103= MEMEnIn2[103:103];
assign MEMRWEnOut2103= MEMRWEnIn2[103:103];
assign MEMAddrOut2103= MEMAddrIn2[623:618];
assign MEMEnOut2104= MEMEnIn2[104:104];
assign MEMRWEnOut2104= MEMRWEnIn2[104:104];
assign MEMAddrOut2104= MEMAddrIn2[629:624];
assign MEMEnOut2105= MEMEnIn2[105:105];
assign MEMRWEnOut2105= MEMRWEnIn2[105:105];
assign MEMAddrOut2105= MEMAddrIn2[635:630];
assign MEMEnOut2106= MEMEnIn2[106:106];
assign MEMRWEnOut2106= MEMRWEnIn2[106:106];
assign MEMAddrOut2106= MEMAddrIn2[641:636];
assign MEMEnOut2107= MEMEnIn2[107:107];
assign MEMRWEnOut2107= MEMRWEnIn2[107:107];
assign MEMAddrOut2107= MEMAddrIn2[647:642];
assign IMEMEnOut2 = IMEMEnIn2;
assign IMEMRWEnOut2 = IMEMRWEnIn2;
assign IMEMAddrOut2 = IMEMAddrIn2;
endmodule
module ArrayTop(
clk,
rst,
dataOut,
dataIn,
configIn,
controlIn,
gControlIn
);
input  clk, rst; 
output [287:0] dataOut; 
input [3455:0] dataIn; 
input [2:0] configIn; 
input [35:0] controlIn; 
input [125:0] gControlIn; 
wire [287:0] topOutputData_w; 
wire [3455:0] topInputData_w; 
wire [2:0] oConfig_w; 
wire [35:0] oControl_w; 
wire [125:0] gControl_w; 
assign dataOut = topOutputData_w; 
assign topInputData_w = dataIn; 
assign oConfig_w = configIn; 
assign oControl_w = controlIn; 
assign gControl_w = gControlIn; 
wire [2:0]MS_OConfigS0_w0;
wire [2:0]MS_IConfigS0_w0;
HA_Reg MS_ConfigS0_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w0),
.DataOut_1(MS_OConfigS0_w0)
);
defparam MS_ConfigS0_0.DataIn_1_BW = 3;
defparam MS_ConfigS0_0.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w0;
wire [3:0]MS_OEnS0_w0;
HA_Reg MS_EnS0_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w0),
.DataOut_1(MS_OEnS0_w0)
);
defparam MS_EnS0_0.DataIn_1_BW = 4;
defparam MS_EnS0_0.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w1;
wire [2:0]MS_IConfigS0_w1;
HA_Reg MS_ConfigS0_1(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w1),
.DataOut_1(MS_OConfigS0_w1)
);
defparam MS_ConfigS0_1.DataIn_1_BW = 3;
defparam MS_ConfigS0_1.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w1;
wire [3:0]MS_OEnS0_w1;
HA_Reg MS_EnS0_1(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w1),
.DataOut_1(MS_OEnS0_w1)
);
defparam MS_EnS0_1.DataIn_1_BW = 4;
defparam MS_EnS0_1.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w2;
wire [2:0]MS_IConfigS0_w2;
HA_Reg MS_ConfigS0_2(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w2),
.DataOut_1(MS_OConfigS0_w2)
);
defparam MS_ConfigS0_2.DataIn_1_BW = 3;
defparam MS_ConfigS0_2.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w2;
wire [3:0]MS_OEnS0_w2;
HA_Reg MS_EnS0_2(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w2),
.DataOut_1(MS_OEnS0_w2)
);
defparam MS_EnS0_2.DataIn_1_BW = 4;
defparam MS_EnS0_2.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w3;
wire [2:0]MS_IConfigS0_w3;
HA_Reg MS_ConfigS0_3(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w3),
.DataOut_1(MS_OConfigS0_w3)
);
defparam MS_ConfigS0_3.DataIn_1_BW = 3;
defparam MS_ConfigS0_3.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w3;
wire [3:0]MS_OEnS0_w3;
HA_Reg MS_EnS0_3(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w3),
.DataOut_1(MS_OEnS0_w3)
);
defparam MS_EnS0_3.DataIn_1_BW = 4;
defparam MS_EnS0_3.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w4;
wire [2:0]MS_IConfigS0_w4;
HA_Reg MS_ConfigS0_4(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w4),
.DataOut_1(MS_OConfigS0_w4)
);
defparam MS_ConfigS0_4.DataIn_1_BW = 3;
defparam MS_ConfigS0_4.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w4;
wire [3:0]MS_OEnS0_w4;
HA_Reg MS_EnS0_4(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w4),
.DataOut_1(MS_OEnS0_w4)
);
defparam MS_EnS0_4.DataIn_1_BW = 4;
defparam MS_EnS0_4.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w5;
wire [2:0]MS_IConfigS0_w5;
HA_Reg MS_ConfigS0_5(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w5),
.DataOut_1(MS_OConfigS0_w5)
);
defparam MS_ConfigS0_5.DataIn_1_BW = 3;
defparam MS_ConfigS0_5.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w5;
wire [3:0]MS_OEnS0_w5;
HA_Reg MS_EnS0_5(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w5),
.DataOut_1(MS_OEnS0_w5)
);
defparam MS_EnS0_5.DataIn_1_BW = 4;
defparam MS_EnS0_5.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w6;
wire [2:0]MS_IConfigS0_w6;
HA_Reg MS_ConfigS0_6(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w6),
.DataOut_1(MS_OConfigS0_w6)
);
defparam MS_ConfigS0_6.DataIn_1_BW = 3;
defparam MS_ConfigS0_6.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w6;
wire [3:0]MS_OEnS0_w6;
HA_Reg MS_EnS0_6(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w6),
.DataOut_1(MS_OEnS0_w6)
);
defparam MS_EnS0_6.DataIn_1_BW = 4;
defparam MS_EnS0_6.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w7;
wire [2:0]MS_IConfigS0_w7;
HA_Reg MS_ConfigS0_7(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w7),
.DataOut_1(MS_OConfigS0_w7)
);
defparam MS_ConfigS0_7.DataIn_1_BW = 3;
defparam MS_ConfigS0_7.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w7;
wire [3:0]MS_OEnS0_w7;
HA_Reg MS_EnS0_7(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w7),
.DataOut_1(MS_OEnS0_w7)
);
defparam MS_EnS0_7.DataIn_1_BW = 4;
defparam MS_EnS0_7.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS0_w8;
wire [2:0]MS_IConfigS0_w8;
HA_Reg MS_ConfigS0_8(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS0_w8),
.DataOut_1(MS_OConfigS0_w8)
);
defparam MS_ConfigS0_8.DataIn_1_BW = 3;
defparam MS_ConfigS0_8.DataOut_1_BW = 3;
wire [3:0]MS_IEnS0_w8;
wire [3:0]MS_OEnS0_w8;
HA_Reg MS_EnS0_8(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS0_w8),
.DataOut_1(MS_OEnS0_w8)
);
defparam MS_EnS0_8.DataIn_1_BW = 4;
defparam MS_EnS0_8.DataOut_1_BW = 4;
wire [2:0]MS_OConfigS1_w0;
wire [2:0]MS_IConfigS1_w0;
HA_Reg MS_ConfigS1_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS1_w0),
.DataOut_1(MS_OConfigS1_w0)
);
defparam MS_ConfigS1_0.DataIn_1_BW = 3;
defparam MS_ConfigS1_0.DataOut_1_BW = 3;
wire [15:0]MS_IEnS1_w0;
wire [15:0]MS_OEnS1_w0;
HA_Reg MS_EnS1_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS1_w0),
.DataOut_1(MS_OEnS1_w0)
);
defparam MS_EnS1_0.DataIn_1_BW = 16;
defparam MS_EnS1_0.DataOut_1_BW = 16;
assign MS_IConfigS0_w0 = MS_OConfigS1_w0;
assign MS_IEnS0_w0 = MS_OEnS1_w0[15:12];
assign MS_IConfigS0_w1 = MS_OConfigS1_w0;
assign MS_IEnS0_w1 = MS_OEnS1_w0[11:8];
assign MS_IConfigS0_w2 = MS_OConfigS1_w0;
assign MS_IEnS0_w2 = MS_OEnS1_w0[7:4];
assign MS_IConfigS0_w3 = MS_OConfigS1_w0;
assign MS_IEnS0_w3 = MS_OEnS1_w0[3:0];
wire [2:0]MS_OConfigS1_w1;
wire [2:0]MS_IConfigS1_w1;
HA_Reg MS_ConfigS1_1(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS1_w1),
.DataOut_1(MS_OConfigS1_w1)
);
defparam MS_ConfigS1_1.DataIn_1_BW = 3;
defparam MS_ConfigS1_1.DataOut_1_BW = 3;
wire [15:0]MS_IEnS1_w1;
wire [15:0]MS_OEnS1_w1;
HA_Reg MS_EnS1_1(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS1_w1),
.DataOut_1(MS_OEnS1_w1)
);
defparam MS_EnS1_1.DataIn_1_BW = 16;
defparam MS_EnS1_1.DataOut_1_BW = 16;
assign MS_IConfigS0_w4 = MS_OConfigS1_w1;
assign MS_IEnS0_w4 = MS_OEnS1_w1[15:12];
assign MS_IConfigS0_w5 = MS_OConfigS1_w1;
assign MS_IEnS0_w5 = MS_OEnS1_w1[11:8];
assign MS_IConfigS0_w6 = MS_OConfigS1_w1;
assign MS_IEnS0_w6 = MS_OEnS1_w1[7:4];
assign MS_IConfigS0_w7 = MS_OConfigS1_w1;
assign MS_IEnS0_w7 = MS_OEnS1_w1[3:0];
wire [2:0]MS_OConfigS1_w2;
wire [2:0]MS_IConfigS1_w2;
HA_Reg MS_ConfigS1_2(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS1_w2),
.DataOut_1(MS_OConfigS1_w2)
);
defparam MS_ConfigS1_2.DataIn_1_BW = 3;
defparam MS_ConfigS1_2.DataOut_1_BW = 3;
wire [3:0]MS_IEnS1_w2;
wire [3:0]MS_OEnS1_w2;
HA_Reg MS_EnS1_2(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS1_w2),
.DataOut_1(MS_OEnS1_w2)
);
defparam MS_EnS1_2.DataIn_1_BW = 4;
defparam MS_EnS1_2.DataOut_1_BW = 4;
assign MS_IConfigS0_w8 = MS_OConfigS1_w2;
assign MS_IEnS0_w8 = MS_OEnS1_w2[3:0];
wire [2:0]MS_OConfigS2_w0;
wire [2:0]MS_IConfigS2_w0;
HA_Reg MS_ConfigS2_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IConfigS2_w0),
.DataOut_1(MS_OConfigS2_w0)
);
defparam MS_ConfigS2_0.DataIn_1_BW = 3;
defparam MS_ConfigS2_0.DataOut_1_BW = 3;
wire [35:0]MS_IEnS2_w0;
wire [35:0]MS_OEnS2_w0;
HA_Reg MS_EnS2_0(
.clk(clk),
.rst(rst),
.DataIn_1(MS_IEnS2_w0),
.DataOut_1(MS_OEnS2_w0)
);
defparam MS_EnS2_0.DataIn_1_BW = 36;
defparam MS_EnS2_0.DataOut_1_BW = 36;
assign MS_IConfigS1_w0 = MS_OConfigS2_w0;
assign MS_IEnS1_w0 = MS_OEnS2_w0[35:20];
assign MS_IConfigS1_w1 = MS_OConfigS2_w0;
assign MS_IEnS1_w1 = MS_OEnS2_w0[19:4];
assign MS_IConfigS1_w2 = MS_OConfigS2_w0;
assign MS_IEnS1_w2 = MS_OEnS2_w0[3:0];
assign MS_IConfigS2_w0 = oConfig_w[2:0]; 
assign MS_IEnS2_w0 = oControl_w;
wire [31:0] V0_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_0_VSTop_Config_Reg_EN; 
wire [2:0] V0_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_0_VSTop_Config_Reg_EN; 
wire [2:0] V1_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_0_VSTop_Config_Reg_EN; 
wire [2:0] V2_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_0_VSTop_Config_Reg_EN; 
wire [2:0] V3_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_0_VSTop_Config_Reg_EN; 
wire [2:0] V4_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_0_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_0_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_0_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_0_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_0_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_0_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_0_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_0_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_0_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_0_VSTop_Config_Reg_EN; 
wire [2:0] V5_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_0_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_0_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_0_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_0_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_0_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_0_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_0_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_0_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_0_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_0_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_0_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V0_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_1_VSTop_Config_Reg_EN; 
wire [2:0] V0_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_1_VSTop_Config_Reg_EN; 
wire [2:0] V1_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_1_VSTop_Config_Reg_EN; 
wire [2:0] V2_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_1_VSTop_Config_Reg_EN; 
wire [2:0] V3_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_1_VSTop_Config_Reg_EN; 
wire [2:0] V4_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_1_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_1_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_1_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_1_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_1_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_1_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_1_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_1_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_1_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_1_VSTop_Config_Reg_EN; 
wire [2:0] V5_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_1_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_1_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_1_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_1_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_1_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_1_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_1_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_1_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_1_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_1_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_1_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V0_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_2_VSTop_Config_Reg_EN; 
wire [2:0] V0_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_2_VSTop_Config_Reg_EN; 
wire [2:0] V1_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_2_VSTop_Config_Reg_EN; 
wire [2:0] V2_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_2_VSTop_Config_Reg_EN; 
wire [2:0] V3_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_2_VSTop_Config_Reg_EN; 
wire [2:0] V4_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_2_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_2_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_2_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_2_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_2_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_2_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_2_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_2_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_2_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_2_VSTop_Config_Reg_EN; 
wire [2:0] V5_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_2_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_2_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_2_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_2_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_2_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_2_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_2_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_2_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_2_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_2_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_2_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V0_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_3_VSTop_Config_Reg_EN; 
wire [2:0] V0_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_3_VSTop_Config_Reg_EN; 
wire [2:0] V1_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_3_VSTop_Config_Reg_EN; 
wire [2:0] V2_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_3_VSTop_Config_Reg_EN; 
wire [2:0] V3_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_3_VSTop_Config_Reg_EN; 
wire [2:0] V4_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_3_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_3_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_3_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_3_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_3_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_3_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_3_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_3_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_3_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_3_VSTop_Config_Reg_EN; 
wire [2:0] V5_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_3_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_3_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_3_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_3_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_3_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_3_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_3_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_3_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_3_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_3_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_3_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V0_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_4_VSTop_Config_Reg_EN; 
wire [2:0] V0_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_4_VSTop_Config_Reg_EN; 
wire [2:0] V1_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_4_VSTop_Config_Reg_EN; 
wire [2:0] V2_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_4_VSTop_Config_Reg_EN; 
wire [2:0] V3_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_4_VSTop_Config_Reg_EN; 
wire [2:0] V4_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_4_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_4_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_4_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_4_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_4_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_4_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_4_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_4_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_4_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_4_VSTop_Config_Reg_EN; 
wire [2:0] V5_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_4_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_4_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_4_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_4_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_4_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_4_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_4_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_4_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_4_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_4_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_4_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V0_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V0_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V0_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V0_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V0_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V0_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V0_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V0_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V0_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V0_5_VSTop_Config_Reg_EN; 
wire [2:0] V0_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V0_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V0_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V0_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V0_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V0_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V0_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V0_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V0_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V0_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V0_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V0_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V0_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V1_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V1_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V1_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V1_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V1_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V1_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V1_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V1_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V1_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V1_5_VSTop_Config_Reg_EN; 
wire [2:0] V1_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V1_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V1_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V1_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V1_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V1_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V1_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V1_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V1_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V1_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V1_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V1_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V1_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V2_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V2_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V2_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V2_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V2_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V2_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V2_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V2_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V2_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V2_5_VSTop_Config_Reg_EN; 
wire [2:0] V2_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V2_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V2_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V2_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V2_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V2_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V2_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V2_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V2_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V2_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V2_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V2_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V2_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V3_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V3_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V3_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V3_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V3_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V3_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V3_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V3_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V3_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V3_5_VSTop_Config_Reg_EN; 
wire [2:0] V3_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V3_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V3_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V3_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V3_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V3_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V3_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V3_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V3_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V3_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V3_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V3_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V3_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V4_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V4_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V4_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V4_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V4_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V4_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V4_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V4_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V4_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V4_5_VSTop_Config_Reg_EN; 
wire [2:0] V4_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V4_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V4_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V4_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V4_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V4_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V4_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V4_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V4_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V4_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V4_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V4_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V4_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

wire [31:0] V5_5_VSTop_VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] V5_5_VSTop_DSE_Solution_L0_GlobalIn0; 
wire [31:0] V5_5_VSTop_DSE_Solution_L0_GlobalIn1; 
wire [31:0] V5_5_VSTop_DSE_Solution_L0_GlobalIn2; 
wire [31:0] V5_5_VSTop_VS_DSE_Solution_L2_t3_O0_3; 
wire [31:0] V5_5_VSTop_VS_DSE_Solution_L5_t5_O0_3; 
wire [0:0] V5_5_VSTop_DSE_Solution_L0_GlobalSel0; 
wire [0:0] V5_5_VSTop_DSE_Solution_L0_GlobalSel1; 
wire [0:0] V5_5_VSTop_DSE_Solution_L0_GlobalSel2; 
wire [0:0] V5_5_VSTop_Config_Reg_EN; 
wire [2:0] V5_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
VSTop V5_5_VSTop( 
.clk(clk),
.rst(rst),
.VSTop_VS_DSE_Solution_L1_t1_In0_1(V5_5_VSTop_VS_DSE_Solution_L1_t1_In0_1),
.VSTop_DSE_Solution_L0_GlobalIn0(V5_5_VSTop_DSE_Solution_L0_GlobalIn0),
.VSTop_DSE_Solution_L0_GlobalIn1(V5_5_VSTop_DSE_Solution_L0_GlobalIn1),
.VSTop_DSE_Solution_L0_GlobalIn2(V5_5_VSTop_DSE_Solution_L0_GlobalIn2),
.VSTop_VS_DSE_Solution_L2_t3_O0_3(V5_5_VSTop_VS_DSE_Solution_L2_t3_O0_3),
.VSTop_VS_DSE_Solution_L5_t5_O0_3(V5_5_VSTop_VS_DSE_Solution_L5_t5_O0_3),
.VSTop_Config_Reg_EN(V5_5_VSTop_Config_Reg_EN),
.VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn(V5_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn),
.VSTop_DSE_Solution_L0_GlobalSel0(V5_5_VSTop_DSE_Solution_L0_GlobalSel0),
.VSTop_DSE_Solution_L0_GlobalSel1(V5_5_VSTop_DSE_Solution_L0_GlobalSel1),
.VSTop_DSE_Solution_L0_GlobalSel2(V5_5_VSTop_DSE_Solution_L0_GlobalSel2)
); 

assign V0_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V0_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V0_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V1_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V1_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V1_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V2_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V2_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V2_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V3_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V3_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V3_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V4_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V4_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V4_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V5_0_VSTop_VS_DSE_Solution_L1_t1_In0_1 = 0;
assign V5_1_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V5_0_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V0_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V0_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V1_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V1_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V2_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V2_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V3_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V3_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V4_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V4_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V5_2_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V5_1_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V0_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V0_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V1_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V1_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V2_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V2_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V3_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V3_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V4_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V4_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V5_3_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V5_2_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V0_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V0_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V1_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V1_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V2_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V2_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V3_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V3_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V4_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V4_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V5_4_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V5_3_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V0_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V0_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V1_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V1_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V2_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V2_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V3_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V3_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V4_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V4_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;
assign V5_5_VSTop_VS_DSE_Solution_L1_t1_In0_1 = V5_4_VSTop_VS_DSE_Solution_L2_t3_O0_3;


assign V0_0_VSTop_Config_Reg_EN = MS_OEnS0_w0[3:3];
assign V0_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w0[2:0];
assign V1_0_VSTop_Config_Reg_EN = MS_OEnS0_w0[2:2];
assign V1_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w0[2:0];
assign V2_0_VSTop_Config_Reg_EN = MS_OEnS0_w0[1:1];
assign V2_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w0[2:0];
assign V3_0_VSTop_Config_Reg_EN = MS_OEnS0_w0[0:0];
assign V3_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w0[2:0];
assign V4_0_VSTop_Config_Reg_EN = MS_OEnS0_w1[3:3];
assign V4_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w1[2:0];
assign V5_0_VSTop_Config_Reg_EN = MS_OEnS0_w1[2:2];
assign V5_0_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w1[2:0];
assign V0_1_VSTop_Config_Reg_EN = MS_OEnS0_w1[1:1];
assign V0_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w1[2:0];
assign V1_1_VSTop_Config_Reg_EN = MS_OEnS0_w1[0:0];
assign V1_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w1[2:0];
assign V2_1_VSTop_Config_Reg_EN = MS_OEnS0_w2[3:3];
assign V2_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w2[2:0];
assign V3_1_VSTop_Config_Reg_EN = MS_OEnS0_w2[2:2];
assign V3_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w2[2:0];
assign V4_1_VSTop_Config_Reg_EN = MS_OEnS0_w2[1:1];
assign V4_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w2[2:0];
assign V5_1_VSTop_Config_Reg_EN = MS_OEnS0_w2[0:0];
assign V5_1_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w2[2:0];
assign V0_2_VSTop_Config_Reg_EN = MS_OEnS0_w3[3:3];
assign V0_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w3[2:0];
assign V1_2_VSTop_Config_Reg_EN = MS_OEnS0_w3[2:2];
assign V1_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w3[2:0];
assign V2_2_VSTop_Config_Reg_EN = MS_OEnS0_w3[1:1];
assign V2_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w3[2:0];
assign V3_2_VSTop_Config_Reg_EN = MS_OEnS0_w3[0:0];
assign V3_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w3[2:0];
assign V4_2_VSTop_Config_Reg_EN = MS_OEnS0_w4[3:3];
assign V4_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w4[2:0];
assign V5_2_VSTop_Config_Reg_EN = MS_OEnS0_w4[2:2];
assign V5_2_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w4[2:0];
assign V0_3_VSTop_Config_Reg_EN = MS_OEnS0_w4[1:1];
assign V0_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w4[2:0];
assign V1_3_VSTop_Config_Reg_EN = MS_OEnS0_w4[0:0];
assign V1_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w4[2:0];
assign V2_3_VSTop_Config_Reg_EN = MS_OEnS0_w5[3:3];
assign V2_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w5[2:0];
assign V3_3_VSTop_Config_Reg_EN = MS_OEnS0_w5[2:2];
assign V3_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w5[2:0];
assign V4_3_VSTop_Config_Reg_EN = MS_OEnS0_w5[1:1];
assign V4_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w5[2:0];
assign V5_3_VSTop_Config_Reg_EN = MS_OEnS0_w5[0:0];
assign V5_3_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w5[2:0];
assign V0_4_VSTop_Config_Reg_EN = MS_OEnS0_w6[3:3];
assign V0_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w6[2:0];
assign V1_4_VSTop_Config_Reg_EN = MS_OEnS0_w6[2:2];
assign V1_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w6[2:0];
assign V2_4_VSTop_Config_Reg_EN = MS_OEnS0_w6[1:1];
assign V2_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w6[2:0];
assign V3_4_VSTop_Config_Reg_EN = MS_OEnS0_w6[0:0];
assign V3_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w6[2:0];
assign V4_4_VSTop_Config_Reg_EN = MS_OEnS0_w7[3:3];
assign V4_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w7[2:0];
assign V5_4_VSTop_Config_Reg_EN = MS_OEnS0_w7[2:2];
assign V5_4_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w7[2:0];
assign V0_5_VSTop_Config_Reg_EN = MS_OEnS0_w7[1:1];
assign V0_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w7[2:0];
assign V1_5_VSTop_Config_Reg_EN = MS_OEnS0_w7[0:0];
assign V1_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w7[2:0];
assign V2_5_VSTop_Config_Reg_EN = MS_OEnS0_w8[3:3];
assign V2_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w8[2:0];
assign V3_5_VSTop_Config_Reg_EN = MS_OEnS0_w8[2:2];
assign V3_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w8[2:0];
assign V4_5_VSTop_Config_Reg_EN = MS_OEnS0_w8[1:1];
assign V4_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w8[2:0];
assign V5_5_VSTop_Config_Reg_EN = MS_OEnS0_w8[0:0];
assign V5_5_VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn = MS_OConfigS0_w8[2:0];
wire [31:0] GIN_0_0_0_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_0_0_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[0:0];
assign GIN_0_0_0_0 = topInputData_w[31:0];
wire [31:0] GIN_0_0_1_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_0_1_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[1:1];
assign GIN_0_0_1_0 = topInputData_w[63:32];
wire [31:0] GIN_0_0_2_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_0_2_0;
assign V0_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[2:2];
assign GIN_0_0_2_0 = topInputData_w[95:64];
wire [31:0] GIN_0_1_0_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_1_0_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[3:3];
assign GIN_0_1_0_0 = topInputData_w[127:96];
wire [31:0] GIN_0_1_1_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_1_1_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[4:4];
assign GIN_0_1_1_0 = topInputData_w[159:128];
wire [31:0] GIN_0_1_2_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_1_2_0;
assign V1_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[5:5];
assign GIN_0_1_2_0 = topInputData_w[191:160];
wire [31:0] GIN_0_2_0_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_2_0_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[6:6];
assign GIN_0_2_0_0 = topInputData_w[223:192];
wire [31:0] GIN_0_2_1_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_2_1_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[7:7];
assign GIN_0_2_1_0 = topInputData_w[255:224];
wire [31:0] GIN_0_2_2_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_2_2_0;
assign V2_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[8:8];
assign GIN_0_2_2_0 = topInputData_w[287:256];
wire [31:0] GIN_0_3_0_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_3_0_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[9:9];
assign GIN_0_3_0_0 = topInputData_w[319:288];
wire [31:0] GIN_0_3_1_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_3_1_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[10:10];
assign GIN_0_3_1_0 = topInputData_w[351:320];
wire [31:0] GIN_0_3_2_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_3_2_0;
assign V3_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[11:11];
assign GIN_0_3_2_0 = topInputData_w[383:352];
wire [31:0] GIN_0_4_0_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_4_0_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[12:12];
assign GIN_0_4_0_0 = topInputData_w[415:384];
wire [31:0] GIN_0_4_1_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_4_1_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[13:13];
assign GIN_0_4_1_0 = topInputData_w[447:416];
wire [31:0] GIN_0_4_2_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_4_2_0;
assign V4_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[14:14];
assign GIN_0_4_2_0 = topInputData_w[479:448];
wire [31:0] GIN_0_5_0_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_0_5_0_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[15:15];
assign GIN_0_5_0_0 = topInputData_w[511:480];
wire [31:0] GIN_0_5_1_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_0_5_1_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[16:16];
assign GIN_0_5_1_0 = topInputData_w[543:512];
wire [31:0] GIN_0_5_2_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_0_5_2_0;
assign V5_0_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[17:17];
assign GIN_0_5_2_0 = topInputData_w[575:544];
wire [31:0] GIN_1_0_0_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_0_0_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[18:18];
assign GIN_1_0_0_0 = topInputData_w[607:576];
wire [31:0] GIN_1_0_1_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_0_1_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[19:19];
assign GIN_1_0_1_0 = topInputData_w[639:608];
wire [31:0] GIN_1_0_2_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_0_2_0;
assign V0_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[20:20];
assign GIN_1_0_2_0 = topInputData_w[671:640];
wire [31:0] GIN_1_1_0_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_1_0_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[21:21];
assign GIN_1_1_0_0 = topInputData_w[703:672];
wire [31:0] GIN_1_1_1_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_1_1_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[22:22];
assign GIN_1_1_1_0 = topInputData_w[735:704];
wire [31:0] GIN_1_1_2_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_1_2_0;
assign V1_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[23:23];
assign GIN_1_1_2_0 = topInputData_w[767:736];
wire [31:0] GIN_1_2_0_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_2_0_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[24:24];
assign GIN_1_2_0_0 = topInputData_w[799:768];
wire [31:0] GIN_1_2_1_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_2_1_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[25:25];
assign GIN_1_2_1_0 = topInputData_w[831:800];
wire [31:0] GIN_1_2_2_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_2_2_0;
assign V2_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[26:26];
assign GIN_1_2_2_0 = topInputData_w[863:832];
wire [31:0] GIN_1_3_0_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_3_0_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[27:27];
assign GIN_1_3_0_0 = topInputData_w[895:864];
wire [31:0] GIN_1_3_1_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_3_1_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[28:28];
assign GIN_1_3_1_0 = topInputData_w[927:896];
wire [31:0] GIN_1_3_2_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_3_2_0;
assign V3_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[29:29];
assign GIN_1_3_2_0 = topInputData_w[959:928];
wire [31:0] GIN_1_4_0_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_4_0_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[30:30];
assign GIN_1_4_0_0 = topInputData_w[991:960];
wire [31:0] GIN_1_4_1_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_4_1_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[31:31];
assign GIN_1_4_1_0 = topInputData_w[1023:992];
wire [31:0] GIN_1_4_2_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_4_2_0;
assign V4_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[32:32];
assign GIN_1_4_2_0 = topInputData_w[1055:1024];
wire [31:0] GIN_1_5_0_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_1_5_0_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[33:33];
assign GIN_1_5_0_0 = topInputData_w[1087:1056];
wire [31:0] GIN_1_5_1_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_1_5_1_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[34:34];
assign GIN_1_5_1_0 = topInputData_w[1119:1088];
wire [31:0] GIN_1_5_2_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_1_5_2_0;
assign V5_1_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[35:35];
assign GIN_1_5_2_0 = topInputData_w[1151:1120];
wire [31:0] GIN_2_0_0_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_0_0_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[36:36];
assign GIN_2_0_0_0 = topInputData_w[1183:1152];
wire [31:0] GIN_2_0_1_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_0_1_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[37:37];
assign GIN_2_0_1_0 = topInputData_w[1215:1184];
wire [31:0] GIN_2_0_2_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_0_2_0;
assign V0_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[38:38];
assign GIN_2_0_2_0 = topInputData_w[1247:1216];
wire [31:0] GIN_2_1_0_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_1_0_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[39:39];
assign GIN_2_1_0_0 = topInputData_w[1279:1248];
wire [31:0] GIN_2_1_1_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_1_1_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[40:40];
assign GIN_2_1_1_0 = topInputData_w[1311:1280];
wire [31:0] GIN_2_1_2_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_1_2_0;
assign V1_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[41:41];
assign GIN_2_1_2_0 = topInputData_w[1343:1312];
wire [31:0] GIN_2_2_0_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_2_0_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[42:42];
assign GIN_2_2_0_0 = topInputData_w[1375:1344];
wire [31:0] GIN_2_2_1_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_2_1_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[43:43];
assign GIN_2_2_1_0 = topInputData_w[1407:1376];
wire [31:0] GIN_2_2_2_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_2_2_0;
assign V2_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[44:44];
assign GIN_2_2_2_0 = topInputData_w[1439:1408];
wire [31:0] GIN_2_3_0_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_3_0_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[45:45];
assign GIN_2_3_0_0 = topInputData_w[1471:1440];
wire [31:0] GIN_2_3_1_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_3_1_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[46:46];
assign GIN_2_3_1_0 = topInputData_w[1503:1472];
wire [31:0] GIN_2_3_2_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_3_2_0;
assign V3_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[47:47];
assign GIN_2_3_2_0 = topInputData_w[1535:1504];
wire [31:0] GIN_2_4_0_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_4_0_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[48:48];
assign GIN_2_4_0_0 = topInputData_w[1567:1536];
wire [31:0] GIN_2_4_1_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_4_1_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[49:49];
assign GIN_2_4_1_0 = topInputData_w[1599:1568];
wire [31:0] GIN_2_4_2_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_4_2_0;
assign V4_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[50:50];
assign GIN_2_4_2_0 = topInputData_w[1631:1600];
wire [31:0] GIN_2_5_0_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_2_5_0_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[51:51];
assign GIN_2_5_0_0 = topInputData_w[1663:1632];
wire [31:0] GIN_2_5_1_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_2_5_1_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[52:52];
assign GIN_2_5_1_0 = topInputData_w[1695:1664];
wire [31:0] GIN_2_5_2_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_2_5_2_0;
assign V5_2_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[53:53];
assign GIN_2_5_2_0 = topInputData_w[1727:1696];
wire [31:0] GIN_3_0_0_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_0_0_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[54:54];
assign GIN_3_0_0_0 = topInputData_w[1759:1728];
wire [31:0] GIN_3_0_1_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_0_1_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[55:55];
assign GIN_3_0_1_0 = topInputData_w[1791:1760];
wire [31:0] GIN_3_0_2_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_0_2_0;
assign V0_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[56:56];
assign GIN_3_0_2_0 = topInputData_w[1823:1792];
wire [31:0] GIN_3_1_0_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_1_0_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[57:57];
assign GIN_3_1_0_0 = topInputData_w[1855:1824];
wire [31:0] GIN_3_1_1_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_1_1_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[58:58];
assign GIN_3_1_1_0 = topInputData_w[1887:1856];
wire [31:0] GIN_3_1_2_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_1_2_0;
assign V1_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[59:59];
assign GIN_3_1_2_0 = topInputData_w[1919:1888];
wire [31:0] GIN_3_2_0_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_2_0_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[60:60];
assign GIN_3_2_0_0 = topInputData_w[1951:1920];
wire [31:0] GIN_3_2_1_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_2_1_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[61:61];
assign GIN_3_2_1_0 = topInputData_w[1983:1952];
wire [31:0] GIN_3_2_2_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_2_2_0;
assign V2_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[62:62];
assign GIN_3_2_2_0 = topInputData_w[2015:1984];
wire [31:0] GIN_3_3_0_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_3_0_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[63:63];
assign GIN_3_3_0_0 = topInputData_w[2047:2016];
wire [31:0] GIN_3_3_1_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_3_1_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[64:64];
assign GIN_3_3_1_0 = topInputData_w[2079:2048];
wire [31:0] GIN_3_3_2_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_3_2_0;
assign V3_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[65:65];
assign GIN_3_3_2_0 = topInputData_w[2111:2080];
wire [31:0] GIN_3_4_0_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_4_0_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[66:66];
assign GIN_3_4_0_0 = topInputData_w[2143:2112];
wire [31:0] GIN_3_4_1_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_4_1_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[67:67];
assign GIN_3_4_1_0 = topInputData_w[2175:2144];
wire [31:0] GIN_3_4_2_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_4_2_0;
assign V4_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[68:68];
assign GIN_3_4_2_0 = topInputData_w[2207:2176];
wire [31:0] GIN_3_5_0_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_3_5_0_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[69:69];
assign GIN_3_5_0_0 = topInputData_w[2239:2208];
wire [31:0] GIN_3_5_1_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_3_5_1_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[70:70];
assign GIN_3_5_1_0 = topInputData_w[2271:2240];
wire [31:0] GIN_3_5_2_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_3_5_2_0;
assign V5_3_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[71:71];
assign GIN_3_5_2_0 = topInputData_w[2303:2272];
wire [31:0] GIN_4_0_0_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_0_0_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[72:72];
assign GIN_4_0_0_0 = topInputData_w[2335:2304];
wire [31:0] GIN_4_0_1_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_0_1_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[73:73];
assign GIN_4_0_1_0 = topInputData_w[2367:2336];
wire [31:0] GIN_4_0_2_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_0_2_0;
assign V0_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[74:74];
assign GIN_4_0_2_0 = topInputData_w[2399:2368];
wire [31:0] GIN_4_1_0_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_1_0_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[75:75];
assign GIN_4_1_0_0 = topInputData_w[2431:2400];
wire [31:0] GIN_4_1_1_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_1_1_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[76:76];
assign GIN_4_1_1_0 = topInputData_w[2463:2432];
wire [31:0] GIN_4_1_2_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_1_2_0;
assign V1_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[77:77];
assign GIN_4_1_2_0 = topInputData_w[2495:2464];
wire [31:0] GIN_4_2_0_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_2_0_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[78:78];
assign GIN_4_2_0_0 = topInputData_w[2527:2496];
wire [31:0] GIN_4_2_1_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_2_1_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[79:79];
assign GIN_4_2_1_0 = topInputData_w[2559:2528];
wire [31:0] GIN_4_2_2_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_2_2_0;
assign V2_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[80:80];
assign GIN_4_2_2_0 = topInputData_w[2591:2560];
wire [31:0] GIN_4_3_0_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_3_0_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[81:81];
assign GIN_4_3_0_0 = topInputData_w[2623:2592];
wire [31:0] GIN_4_3_1_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_3_1_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[82:82];
assign GIN_4_3_1_0 = topInputData_w[2655:2624];
wire [31:0] GIN_4_3_2_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_3_2_0;
assign V3_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[83:83];
assign GIN_4_3_2_0 = topInputData_w[2687:2656];
wire [31:0] GIN_4_4_0_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_4_0_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[84:84];
assign GIN_4_4_0_0 = topInputData_w[2719:2688];
wire [31:0] GIN_4_4_1_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_4_1_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[85:85];
assign GIN_4_4_1_0 = topInputData_w[2751:2720];
wire [31:0] GIN_4_4_2_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_4_2_0;
assign V4_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[86:86];
assign GIN_4_4_2_0 = topInputData_w[2783:2752];
wire [31:0] GIN_4_5_0_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_4_5_0_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[87:87];
assign GIN_4_5_0_0 = topInputData_w[2815:2784];
wire [31:0] GIN_4_5_1_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_4_5_1_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[88:88];
assign GIN_4_5_1_0 = topInputData_w[2847:2816];
wire [31:0] GIN_4_5_2_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_4_5_2_0;
assign V5_4_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[89:89];
assign GIN_4_5_2_0 = topInputData_w[2879:2848];
wire [31:0] GIN_5_0_0_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_0_0_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[90:90];
assign GIN_5_0_0_0 = topInputData_w[2911:2880];
wire [31:0] GIN_5_0_1_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_0_1_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[91:91];
assign GIN_5_0_1_0 = topInputData_w[2943:2912];
wire [31:0] GIN_5_0_2_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_0_2_0;
assign V0_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[92:92];
assign GIN_5_0_2_0 = topInputData_w[2975:2944];
wire [31:0] GIN_5_1_0_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_1_0_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[93:93];
assign GIN_5_1_0_0 = topInputData_w[3007:2976];
wire [31:0] GIN_5_1_1_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_1_1_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[94:94];
assign GIN_5_1_1_0 = topInputData_w[3039:3008];
wire [31:0] GIN_5_1_2_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_1_2_0;
assign V1_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[95:95];
assign GIN_5_1_2_0 = topInputData_w[3071:3040];
wire [31:0] GIN_5_2_0_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_2_0_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[96:96];
assign GIN_5_2_0_0 = topInputData_w[3103:3072];
wire [31:0] GIN_5_2_1_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_2_1_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[97:97];
assign GIN_5_2_1_0 = topInputData_w[3135:3104];
wire [31:0] GIN_5_2_2_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_2_2_0;
assign V2_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[98:98];
assign GIN_5_2_2_0 = topInputData_w[3167:3136];
wire [31:0] GIN_5_3_0_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_3_0_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[99:99];
assign GIN_5_3_0_0 = topInputData_w[3199:3168];
wire [31:0] GIN_5_3_1_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_3_1_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[100:100];
assign GIN_5_3_1_0 = topInputData_w[3231:3200];
wire [31:0] GIN_5_3_2_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_3_2_0;
assign V3_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[101:101];
assign GIN_5_3_2_0 = topInputData_w[3263:3232];
wire [31:0] GIN_5_4_0_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_4_0_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[102:102];
assign GIN_5_4_0_0 = topInputData_w[3295:3264];
wire [31:0] GIN_5_4_1_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_4_1_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[103:103];
assign GIN_5_4_1_0 = topInputData_w[3327:3296];
wire [31:0] GIN_5_4_2_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_4_2_0;
assign V4_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[104:104];
assign GIN_5_4_2_0 = topInputData_w[3359:3328];
wire [31:0] GIN_5_5_0_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalIn0 = GIN_5_5_0_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalSel0 = gControl_w[105:105];
assign GIN_5_5_0_0 = topInputData_w[3391:3360];
wire [31:0] GIN_5_5_1_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalIn1 = GIN_5_5_1_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalSel1 = gControl_w[106:106];
assign GIN_5_5_1_0 = topInputData_w[3423:3392];
wire [31:0] GIN_5_5_2_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalIn2 = GIN_5_5_2_0;
assign V5_5_VSTop_DSE_Solution_L0_GlobalSel2 = gControl_w[107:107];
assign GIN_5_5_2_0 = topInputData_w[3455:3424];
wire [31:0] gRW0_1;
assign gRW0_1 = V0_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW0_2;
assign gRW0_2 = V1_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW0_3;
assign gRW0_3 = V0_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW0_4;
assign gRW0_4 = V1_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut0;
wire [1:0] grSel0;
HA_4IM grC0(
.sel(grSel0),
.DataOut_1(grOut0),
.DataIn_1(gRW0_1),
.DataIn_2(gRW0_2),
.DataIn_3(gRW0_3),
.DataIn_4(gRW0_4)
);
defparam   grC0.Mux_BW = 32;
assign topOutputData_w[31:0] = grOut0;
assign grSel0 = gControl_w[109:108];
wire [31:0] gRW1_1;
assign gRW1_1 = V2_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW1_2;
assign gRW1_2 = V3_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW1_3;
assign gRW1_3 = V2_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW1_4;
assign gRW1_4 = V3_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut1;
wire [1:0] grSel1;
HA_4IM grC1(
.sel(grSel1),
.DataOut_1(grOut1),
.DataIn_1(gRW1_1),
.DataIn_2(gRW1_2),
.DataIn_3(gRW1_3),
.DataIn_4(gRW1_4)
);
defparam   grC1.Mux_BW = 32;
assign topOutputData_w[63:32] = grOut1;
assign grSel1 = gControl_w[111:110];
wire [31:0] gRW2_1;
assign gRW2_1 = V4_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW2_2;
assign gRW2_2 = V5_0_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW2_3;
assign gRW2_3 = V4_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW2_4;
assign gRW2_4 = V5_1_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut2;
wire [1:0] grSel2;
HA_4IM grC2(
.sel(grSel2),
.DataOut_1(grOut2),
.DataIn_1(gRW2_1),
.DataIn_2(gRW2_2),
.DataIn_3(gRW2_3),
.DataIn_4(gRW2_4)
);
defparam   grC2.Mux_BW = 32;
assign topOutputData_w[95:64] = grOut2;
assign grSel2 = gControl_w[113:112];
wire [31:0] gRW3_1;
assign gRW3_1 = V0_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW3_2;
assign gRW3_2 = V1_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW3_3;
assign gRW3_3 = V0_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW3_4;
assign gRW3_4 = V1_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut3;
wire [1:0] grSel3;
HA_4IM grC3(
.sel(grSel3),
.DataOut_1(grOut3),
.DataIn_1(gRW3_1),
.DataIn_2(gRW3_2),
.DataIn_3(gRW3_3),
.DataIn_4(gRW3_4)
);
defparam   grC3.Mux_BW = 32;
assign topOutputData_w[127:96] = grOut3;
assign grSel3 = gControl_w[115:114];
wire [31:0] gRW4_1;
assign gRW4_1 = V2_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW4_2;
assign gRW4_2 = V3_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW4_3;
assign gRW4_3 = V2_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW4_4;
assign gRW4_4 = V3_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut4;
wire [1:0] grSel4;
HA_4IM grC4(
.sel(grSel4),
.DataOut_1(grOut4),
.DataIn_1(gRW4_1),
.DataIn_2(gRW4_2),
.DataIn_3(gRW4_3),
.DataIn_4(gRW4_4)
);
defparam   grC4.Mux_BW = 32;
assign topOutputData_w[159:128] = grOut4;
assign grSel4 = gControl_w[117:116];
wire [31:0] gRW5_1;
assign gRW5_1 = V4_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW5_2;
assign gRW5_2 = V5_2_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW5_3;
assign gRW5_3 = V4_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW5_4;
assign gRW5_4 = V5_3_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut5;
wire [1:0] grSel5;
HA_4IM grC5(
.sel(grSel5),
.DataOut_1(grOut5),
.DataIn_1(gRW5_1),
.DataIn_2(gRW5_2),
.DataIn_3(gRW5_3),
.DataIn_4(gRW5_4)
);
defparam   grC5.Mux_BW = 32;
assign topOutputData_w[191:160] = grOut5;
assign grSel5 = gControl_w[119:118];
wire [31:0] gRW6_1;
assign gRW6_1 = V0_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW6_2;
assign gRW6_2 = V1_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW6_3;
assign gRW6_3 = V0_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW6_4;
assign gRW6_4 = V1_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut6;
wire [1:0] grSel6;
HA_4IM grC6(
.sel(grSel6),
.DataOut_1(grOut6),
.DataIn_1(gRW6_1),
.DataIn_2(gRW6_2),
.DataIn_3(gRW6_3),
.DataIn_4(gRW6_4)
);
defparam   grC6.Mux_BW = 32;
assign topOutputData_w[223:192] = grOut6;
assign grSel6 = gControl_w[121:120];
wire [31:0] gRW7_1;
assign gRW7_1 = V2_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW7_2;
assign gRW7_2 = V3_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW7_3;
assign gRW7_3 = V2_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW7_4;
assign gRW7_4 = V3_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut7;
wire [1:0] grSel7;
HA_4IM grC7(
.sel(grSel7),
.DataOut_1(grOut7),
.DataIn_1(gRW7_1),
.DataIn_2(gRW7_2),
.DataIn_3(gRW7_3),
.DataIn_4(gRW7_4)
);
defparam   grC7.Mux_BW = 32;
assign topOutputData_w[255:224] = grOut7;
assign grSel7 = gControl_w[123:122];
wire [31:0] gRW8_1;
assign gRW8_1 = V4_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW8_2;
assign gRW8_2 = V5_4_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW8_3;
assign gRW8_3 = V4_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] gRW8_4;
assign gRW8_4 = V5_5_VSTop_VS_DSE_Solution_L5_t5_O0_3;
wire [31:0] grOut8;
wire [1:0] grSel8;
HA_4IM grC8(
.sel(grSel8),
.DataOut_1(grOut8),
.DataIn_1(gRW8_1),
.DataIn_2(gRW8_2),
.DataIn_3(gRW8_3),
.DataIn_4(gRW8_4)
);
defparam   grC8.Mux_BW = 32;
assign topOutputData_w[287:256] = grOut8;
assign grSel8 = gControl_w[125:124];
endmodule
module VSTop( 
clk,
rst,
VSTop_VS_DSE_Solution_L1_t1_In0_1,
VSTop_DSE_Solution_L0_GlobalIn0,
VSTop_DSE_Solution_L0_GlobalIn1,
VSTop_DSE_Solution_L0_GlobalIn2,
VSTop_VS_DSE_Solution_L2_t3_O0_3,
VSTop_VS_DSE_Solution_L5_t5_O0_3,
VSTop_Config_Reg_EN,
VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn,
VSTop_DSE_Solution_L0_GlobalSel0,
VSTop_DSE_Solution_L0_GlobalSel1,
VSTop_DSE_Solution_L0_GlobalSel2
); 

input clk;
input rst;
input [31:0] VSTop_DSE_Solution_L0_GlobalIn0; 
input [31:0] VSTop_DSE_Solution_L0_GlobalIn1; 
input [31:0] VSTop_DSE_Solution_L0_GlobalIn2; 
input [31:0] VSTop_VS_DSE_Solution_L1_t1_In0_1; 
output [31:0] VSTop_VS_DSE_Solution_L2_t3_O0_3; 
output [31:0] VSTop_VS_DSE_Solution_L5_t5_O0_3; 
input [0:0] VSTop_DSE_Solution_L0_GlobalSel0; 
input [0:0] VSTop_DSE_Solution_L0_GlobalSel1; 
input [0:0] VSTop_DSE_Solution_L0_GlobalSel2; 
input [0:0] VSTop_Config_Reg_EN; 
input [2:0] VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn; 
wire [31:0] VS_DSE_Solution_L0_n0_HA_IN_1; 
wire [31:0] VS_DSE_Solution_L0_n0_HA_IN_2; 
wire [31:0] VS_DSE_Solution_L0_n0_HA_IN_3; 
wire [31:0] VS_DSE_Solution_L0_GlobalIn0; 
wire [31:0] VS_DSE_Solution_L0_GlobalIn1; 
wire [31:0] VS_DSE_Solution_L0_GlobalIn2; 
wire [31:0] VS_DSE_Solution_L0_n0_HA_OW_4; 
wire [0:0] VS_DSE_Solution_L0_GlobalSel0; 
wire [0:0] VS_DSE_Solution_L0_GlobalSel1; 
wire [0:0] VS_DSE_Solution_L0_GlobalSel2; 
wire [0:0] VS_DSE_Solution_L0_Config_Reg_EN; 
wire [2:0] VS_DSE_Solution_L0_Config_Reg_InstIn; 
DSE_Solution_L0 VS_DSE_Solution_L0( 
.clk(clk),
.rst(rst),
.DSE_Solution_L0_n0_HA_IN_1(VS_DSE_Solution_L0_n0_HA_IN_1),
.DSE_Solution_L0_n0_HA_IN_2(VS_DSE_Solution_L0_n0_HA_IN_2),
.DSE_Solution_L0_n0_HA_IN_3(VS_DSE_Solution_L0_n0_HA_IN_3),
.DSE_Solution_L0_GlobalIn0(VS_DSE_Solution_L0_GlobalIn0),
.DSE_Solution_L0_GlobalIn1(VS_DSE_Solution_L0_GlobalIn1),
.DSE_Solution_L0_GlobalIn2(VS_DSE_Solution_L0_GlobalIn2),
.DSE_Solution_L0_n0_HA_OW_4(VS_DSE_Solution_L0_n0_HA_OW_4),
.DSE_Solution_L0_Config_Reg_EN(VS_DSE_Solution_L0_Config_Reg_EN),
.DSE_Solution_L0_Config_Reg_InstIn(VS_DSE_Solution_L0_Config_Reg_InstIn),
.DSE_Solution_L0_GlobalSel0(VS_DSE_Solution_L0_GlobalSel0),
.DSE_Solution_L0_GlobalSel1(VS_DSE_Solution_L0_GlobalSel1),
.DSE_Solution_L0_GlobalSel2(VS_DSE_Solution_L0_GlobalSel2)
); 

assign VS_DSE_Solution_L0_GlobalIn0 = VSTop_DSE_Solution_L0_GlobalIn0;
assign VS_DSE_Solution_L0_GlobalIn1 = VSTop_DSE_Solution_L0_GlobalIn1;
assign VS_DSE_Solution_L0_GlobalIn2 = VSTop_DSE_Solution_L0_GlobalIn2;
assign VS_DSE_Solution_L0_GlobalSel0 = VSTop_DSE_Solution_L0_GlobalSel0;
assign VS_DSE_Solution_L0_GlobalSel1 = VSTop_DSE_Solution_L0_GlobalSel1;
assign VS_DSE_Solution_L0_GlobalSel2 = VSTop_DSE_Solution_L0_GlobalSel2;
wire [31:0] VS_DSE_Solution_L1_t1_In0_1; 
wire [31:0] VS_DSE_Solution_L1_t5_O0_3; 
wire [31:0] VS_DSE_Solution_L1_t5_O1_4; 
DSE_Solution_L1 VS_DSE_Solution_L1( 
.clk(clk),
.rst(rst),
.DSE_Solution_L1_t1_In0_1(VS_DSE_Solution_L1_t1_In0_1),
.DSE_Solution_L1_t5_O0_3(VS_DSE_Solution_L1_t5_O0_3),
.DSE_Solution_L1_t5_O1_4(VS_DSE_Solution_L1_t5_O1_4)
); 

wire [31:0] VS_DSE_Solution_L2_t5_In0_1; 
wire [31:0] VS_DSE_Solution_L2_t3_O0_3; 
DSE_Solution_L2 VS_DSE_Solution_L2( 
.clk(clk),
.rst(rst),
.DSE_Solution_L2_t5_In0_1(VS_DSE_Solution_L2_t5_In0_1),
.DSE_Solution_L2_t3_O0_3(VS_DSE_Solution_L2_t3_O0_3)
); 

wire [31:0] VS_DSE_Solution_L3_t5_In0_1; 
wire [31:0] VS_DSE_Solution_L3_t5_O0_3; 
DSE_Solution_L3 VS_DSE_Solution_L3( 
.clk(clk),
.rst(rst),
.DSE_Solution_L3_t5_In0_1(VS_DSE_Solution_L3_t5_In0_1),
.DSE_Solution_L3_t5_O0_3(VS_DSE_Solution_L3_t5_O0_3)
); 

wire [31:0] VS_DSE_Solution_L4_t5_In0_1; 
wire [31:0] VS_DSE_Solution_L4_t5_O0_3; 
DSE_Solution_L4 VS_DSE_Solution_L4( 
.clk(clk),
.rst(rst),
.DSE_Solution_L4_t5_In0_1(VS_DSE_Solution_L4_t5_In0_1),
.DSE_Solution_L4_t5_O0_3(VS_DSE_Solution_L4_t5_O0_3)
); 

wire [31:0] VS_DSE_Solution_L5_t5_In0_1; 
wire [31:0] VS_DSE_Solution_L5_t5_O0_3; 
DSE_Solution_L5 VS_DSE_Solution_L5( 
.clk(clk),
.rst(rst),
.DSE_Solution_L5_t5_In0_1(VS_DSE_Solution_L5_t5_In0_1),
.DSE_Solution_L5_t5_O0_3(VS_DSE_Solution_L5_t5_O0_3)
); 

assign VSTop_VS_DSE_Solution_L5_t5_O0_3 = VS_DSE_Solution_L5_t5_O0_3;
assign VS_DSE_Solution_L5_t5_In0_1 = VS_DSE_Solution_L0_n0_HA_OW_4;
assign VS_DSE_Solution_L0_Config_Reg_InstIn = VSTop_VS_DSE_Solution_L0_Config_Reg_InstIn;
assign VS_DSE_Solution_L0_Config_Reg_EN = VSTop_Config_Reg_EN;


assign VS_DSE_Solution_L0_n0_HA_IN_1 = VS_DSE_Solution_L1_t5_O0_3;
assign VS_DSE_Solution_L0_n0_HA_IN_2 = VS_DSE_Solution_L1_t5_O1_4;
assign VS_DSE_Solution_L1_t1_In0_1 = VSTop_VS_DSE_Solution_L1_t1_In0_1;


assign VSTop_VS_DSE_Solution_L2_t3_O0_3 = VS_DSE_Solution_L2_t3_O0_3;


assign VS_DSE_Solution_L2_t5_In0_1 = VS_DSE_Solution_L3_t5_O0_3;


assign VS_DSE_Solution_L3_t5_In0_1 = VS_DSE_Solution_L4_t5_O0_3;


assign VS_DSE_Solution_L4_t5_In0_1 = VS_DSE_Solution_L5_t5_O0_3;


endmodule
module DSE_Solution_L0( 
clk,
rst,
DSE_Solution_L0_n0_HA_IN_1,
DSE_Solution_L0_n0_HA_IN_2,
DSE_Solution_L0_n0_HA_IN_3,
DSE_Solution_L0_GlobalIn0,
DSE_Solution_L0_GlobalIn1,
DSE_Solution_L0_GlobalIn2,
DSE_Solution_L0_n0_HA_OW_4,
DSE_Solution_L0_Config_Reg_EN,
DSE_Solution_L0_Config_Reg_InstIn,
DSE_Solution_L0_GlobalSel0,
DSE_Solution_L0_GlobalSel1,
DSE_Solution_L0_GlobalSel2
); 

input clk;
input rst;
input [31:0] DSE_Solution_L0_GlobalIn0; 
input [31:0] DSE_Solution_L0_GlobalIn1; 
input [31:0] DSE_Solution_L0_GlobalIn2; 
input [31:0] DSE_Solution_L0_n0_HA_IN_1; 
input [31:0] DSE_Solution_L0_n0_HA_IN_2; 
input [31:0] DSE_Solution_L0_n0_HA_IN_3; 
output [31:0] DSE_Solution_L0_n0_HA_OW_4; 
input [0:0] DSE_Solution_L0_GlobalSel0; 
input [0:0] DSE_Solution_L0_GlobalSel1; 
input [0:0] DSE_Solution_L0_GlobalSel2; 
input [0:0] DSE_Solution_L0_Config_Reg_EN; 
input [2:0] DSE_Solution_L0_Config_Reg_InstIn; 
wire [31:0] n0_HA_IN_1_WDataIn_1;
assign n0_HA_IN_1_WDataIn_1 = DSE_Solution_L0_n0_HA_IN_1;
defparam n0_HA_IN_1.DataIn_1_BW = 32;
wire [31:0] n0_HA_IN_1_WDataIn_2;
assign n0_HA_IN_1_WDataIn_2 = DSE_Solution_L0_GlobalIn0;
defparam n0_HA_IN_1.DataIn_2_BW = 32;
wire [31:0] n0_HA_IN_1_WDataOut_1;
defparam n0_HA_IN_1.DataOut_1_BW = 32;
assign n0_HA_IN_1_Wsel = DSE_Solution_L0_GlobalSel0;
CADA_IN n0_HA_IN_1 (
	.clk( clk ) ,
	.rst( rst ) ,
	.DataIn_1(n0_HA_IN_1_WDataIn_1) ,
	.DataIn_2(n0_HA_IN_1_WDataIn_2) ,
	.DataOut_1(n0_HA_IN_1_WDataOut_1) ,
	.sel(n0_HA_IN_1_Wsel) 
);
wire [31:0] n0_HA_IN_2_WDataIn_1;
assign n0_HA_IN_2_WDataIn_1 = DSE_Solution_L0_n0_HA_IN_2;
defparam n0_HA_IN_2.DataIn_1_BW = 32;
wire [31:0] n0_HA_IN_2_WDataIn_2;
assign n0_HA_IN_2_WDataIn_2 = DSE_Solution_L0_GlobalIn1;
defparam n0_HA_IN_2.DataIn_2_BW = 32;
wire [31:0] n0_HA_IN_2_WDataOut_1;
defparam n0_HA_IN_2.DataOut_1_BW = 32;
assign n0_HA_IN_2_Wsel = DSE_Solution_L0_GlobalSel1;
CADA_IN n0_HA_IN_2 (
	.clk( clk ) ,
	.rst( rst ) ,
	.DataIn_1(n0_HA_IN_2_WDataIn_1) ,
	.DataIn_2(n0_HA_IN_2_WDataIn_2) ,
	.DataOut_1(n0_HA_IN_2_WDataOut_1) ,
	.sel(n0_HA_IN_2_Wsel) 
);
wire [31:0] n0_HA_IN_3_WDataIn_1;
assign n0_HA_IN_3_WDataIn_1 = DSE_Solution_L0_n0_HA_IN_3;
defparam n0_HA_IN_3.DataIn_1_BW = 32;
wire [31:0] n0_HA_IN_3_WDataIn_2;
assign n0_HA_IN_3_WDataIn_2 = DSE_Solution_L0_GlobalIn2;
defparam n0_HA_IN_3.DataIn_2_BW = 32;
wire [31:0] n0_HA_IN_3_WDataOut_1;
defparam n0_HA_IN_3.DataOut_1_BW = 32;
assign n0_HA_IN_3_Wsel = DSE_Solution_L0_GlobalSel2;
CADA_IN n0_HA_IN_3 (
	.clk( clk ) ,
	.rst( rst ) ,
	.DataIn_1(n0_HA_IN_3_WDataIn_1) ,
	.DataIn_2(n0_HA_IN_3_WDataIn_2) ,
	.DataOut_1(n0_HA_IN_3_WDataOut_1) ,
	.sel(n0_HA_IN_3_Wsel) 
);
wire [31:0] n0_HA_OW_4_WDataIn_1;
defparam n0_HA_OW_4.DataIn_1_BW = 32;
wire [31:0] n0_HA_OW_4_WDataOut_1;
assign DSE_Solution_L0_n0_HA_OW_4 = n0_HA_OW_4_WDataOut_1;
defparam n0_HA_OW_4.DataOut_1_BW = 32;
HA_OW n0_HA_OW_4 (
	.DataIn_1(n0_HA_OW_4_WDataIn_1) ,
	.DataOut_1(n0_HA_OW_4_WDataOut_1) 
);
wire [31:0] n0_CADA_ADD_5_WDataIn_1;
defparam n0_CADA_ADD_5.DataIn_1_BW = 32;
wire [31:0] n0_CADA_ADD_5_WDataIn_2;
defparam n0_CADA_ADD_5.DataIn_2_BW = 32;
wire [31:0] n0_CADA_ADD_5_WDataOut_1;
wire [31:0] n0_CADA_ADD_5_DataOut_1_latency_1_WDataIn_1;
wire [31:0] n0_CADA_ADD_5_DataOut_1_latency_1_WDataOut_1;
assign n0_CADA_ADD_5_DataOut_1_latency_1_WDataIn_1 = n0_CADA_ADD_5_WDataOut_1;
HA_Reg n0_CADA_ADD_5_DataOut_1_latency_1 (
	.clk( clk ) ,
	.rst( rst ) ,
	.DataIn_1(n0_CADA_ADD_5_DataOut_1_latency_1_WDataIn_1) ,
	.DataOut_1(n0_CADA_ADD_5_DataOut_1_latency_1_WDataOut_1) 
);
defparam n0_CADA_ADD_5_DataOut_1_latency_1.DataIn_1_BW = 32;
defparam n0_CADA_ADD_5_DataOut_1_latency_1.DataOut_1_BW = 32;
defparam n0_CADA_ADD_5.DataOut_1_BW = 32;
CADA_ADD n0_CADA_ADD_5 (
	.DataIn_1(n0_CADA_ADD_5_WDataIn_1) ,
	.DataIn_2(n0_CADA_ADD_5_WDataIn_2) ,
	.DataOut_1(n0_CADA_ADD_5_WDataOut_1) 
);
wire [31:0] n0_CADA_Mult_6_WDataIn_1;
defparam n0_CADA_Mult_6.DataIn_1_BW = 32;
wire [31:0] n0_CADA_Mult_6_WDataIn_2;
defparam n0_CADA_Mult_6.DataIn_2_BW = 32;
wire [31:0] n0_CADA_Mult_6_WDataOut_1;
wire [31:0] n0_CADA_Mult_6_DataOut_1_latency_1_WDataIn_1;
wire [31:0] n0_CADA_Mult_6_DataOut_1_latency_1_WDataOut_1;
assign n0_CADA_Mult_6_DataOut_1_latency_1_WDataIn_1 = n0_CADA_Mult_6_WDataOut_1;
HA_Reg n0_CADA_Mult_6_DataOut_1_latency_1 (
	.clk( clk ) ,
	.rst( rst ) ,
	.DataIn_1(n0_CADA_Mult_6_DataOut_1_latency_1_WDataIn_1) ,
	.DataOut_1(n0_CADA_Mult_6_DataOut_1_latency_1_WDataOut_1) 
);
defparam n0_CADA_Mult_6_DataOut_1_latency_1.DataIn_1_BW = 32;
defparam n0_CADA_Mult_6_DataOut_1_latency_1.DataOut_1_BW = 32;
defparam n0_CADA_Mult_6.DataOut_1_BW = 32;
CADA_Mult n0_CADA_Mult_6 (
	.DataOut_1(n0_CADA_Mult_6_WDataOut_1) ,
	.DataIn_1(n0_CADA_Mult_6_WDataIn_1) ,
	.DataIn_2(n0_CADA_Mult_6_WDataIn_2) 
);
wire [31:0] LogicMux_1_WDataIn_1;
wire [31:0] LogicMux_1_WDataIn_2;
wire [31:0] LogicMux_1_WDataOut_1;
wire [0:0] LogicMux_1_Wsel;
HA_2IM LogicMux_1 (
	.DataIn_1(LogicMux_1_WDataIn_1) ,
	.DataIn_2(LogicMux_1_WDataIn_2) ,
	.DataOut_1(LogicMux_1_WDataOut_1) ,
	.sel(LogicMux_1_Wsel) 
);
defparam LogicMux_1.Mux_BW = 32;
wire [31:0] LogicMux_2_WDataIn_1;
wire [31:0] LogicMux_2_WDataIn_2;
wire [31:0] LogicMux_2_WDataOut_1;
wire [0:0] LogicMux_2_Wsel;
HA_2IM LogicMux_2 (
	.DataIn_1(LogicMux_2_WDataIn_1) ,
	.DataIn_2(LogicMux_2_WDataIn_2) ,
	.DataOut_1(LogicMux_2_WDataOut_1) ,
	.sel(LogicMux_2_Wsel) 
);
defparam LogicMux_2.Mux_BW = 32;
wire [31:0] LogicMux_3_WDataIn_1;
wire [31:0] LogicMux_3_WDataIn_2;
wire [31:0] LogicMux_3_WDataOut_1;
wire [0:0] LogicMux_3_Wsel;
HA_2IM LogicMux_3 (
	.DataIn_1(LogicMux_3_WDataIn_1) ,
	.DataIn_2(LogicMux_3_WDataIn_2) ,
	.DataOut_1(LogicMux_3_WDataOut_1) ,
	.sel(LogicMux_3_Wsel) 
);
defparam LogicMux_3.Mux_BW = 32;

// Connect child module input to parent module output 

assign n0_CADA_Mult_6_WDataIn_1 = n0_HA_IN_1_WDataOut_1;
assign LogicMux_2_WDataIn_1 = n0_HA_IN_2_WDataOut_1;
assign n0_CADA_ADD_5_WDataIn_1 = LogicMux_2_WDataOut_1;
assign LogicMux_3_WDataIn_1 = n0_HA_IN_2_WDataOut_1;
assign n0_CADA_Mult_6_WDataIn_2 = LogicMux_3_WDataOut_1;

// Connect child module input to parent module output 

assign n0_CADA_ADD_5_WDataIn_2 = n0_HA_IN_3_WDataOut_1;
assign LogicMux_1_WDataIn_1 = n0_CADA_ADD_5_DataOut_1_latency_1_WDataOut_1;
assign n0_HA_OW_4_WDataIn_1 = LogicMux_1_WDataOut_1;
assign LogicMux_3_WDataIn_2 = n0_CADA_ADD_5_DataOut_1_latency_1_WDataOut_1;
assign LogicMux_1_WDataIn_2 = n0_CADA_Mult_6_DataOut_1_latency_1_WDataOut_1;
assign LogicMux_2_WDataIn_2 = n0_CADA_Mult_6_DataOut_1_latency_1_WDataOut_1;
wire [2:0] Config_Reg_WInstOut;
wire [2:0] Config_Reg_WInstIn;
wire [0:0] Config_Reg_WEN;
assign LogicMux_1_Wsel = Config_Reg_WInstOut[0:0]; 
assign LogicMux_2_Wsel = Config_Reg_WInstOut[1:1]; 
assign LogicMux_3_Wsel = Config_Reg_WInstOut[2:2]; 
HA_CReg Config_Reg (
	.clk( clk ) ,
	.rst( rst ) ,
	.InstIn(Config_Reg_WInstIn) ,
	.InstOut(Config_Reg_WInstOut) ,
	.EN(Config_Reg_WEN) 
);
defparam Config_Reg.Inst_BW = 3;
assign Config_Reg_WEN = DSE_Solution_L0_Config_Reg_EN;
assign Config_Reg_WInstIn = DSE_Solution_L0_Config_Reg_InstIn;
endmodule

module DSE_Solution_L1( 
clk,
rst,
DSE_Solution_L1_t1_In0_1,
DSE_Solution_L1_t5_O0_3,
DSE_Solution_L1_t5_O1_4
); 

input clk;
input rst;
input [31:0] DSE_Solution_L1_t1_In0_1; 
output [31:0] DSE_Solution_L1_t5_O0_3; 
output [31:0] DSE_Solution_L1_t5_O1_4; 
wire [31:0] t1_In0_1_WDataIn_1;
assign t1_In0_1_WDataIn_1 = DSE_Solution_L1_t1_In0_1;
defparam t1_In0_1.DataIn_1_BW = 32;
wire [31:0] t1_In0_1_WDataOut_1;
defparam t1_In0_1.DataOut_1_BW = 32;
HA_INW t1_In0_1 (
	.DataIn_1(t1_In0_1_WDataIn_1) ,
	.DataOut_1(t1_In0_1_WDataOut_1) 
);
wire [31:0] Token0_2_WDataIn_1;
defparam Token0_2.DataIn_1_BW = 32;
wire [31:0] Token0_2_WDataOut_1;
defparam Token0_2.DataOut_1_BW = 32;
HA_TW Token0_2 (
	.DataIn_1(Token0_2_WDataIn_1) ,
	.DataOut_1(Token0_2_WDataOut_1) 
);
wire [31:0] t5_O0_3_WDataIn_1;
defparam t5_O0_3.DataIn_1_BW = 32;
wire [31:0] t5_O0_3_WDataOut_1;
assign DSE_Solution_L1_t5_O0_3 = t5_O0_3_WDataOut_1;
defparam t5_O0_3.DataOut_1_BW = 32;
HA_OW t5_O0_3 (
	.DataIn_1(t5_O0_3_WDataIn_1) ,
	.DataOut_1(t5_O0_3_WDataOut_1) 
);
wire [31:0] t5_O1_4_WDataIn_1;
defparam t5_O1_4.DataIn_1_BW = 32;
wire [31:0] t5_O1_4_WDataOut_1;
assign DSE_Solution_L1_t5_O1_4 = t5_O1_4_WDataOut_1;
defparam t5_O1_4.DataOut_1_BW = 32;
HA_OW t5_O1_4 (
	.DataIn_1(t5_O1_4_WDataIn_1) ,
	.DataOut_1(t5_O1_4_WDataOut_1) 
);

// Connect child module input to parent module output 

assign Token0_2_WDataIn_1 = t1_In0_1_WDataOut_1;

// Connect child module input to parent module output 

assign t5_O0_3_WDataIn_1 = Token0_2_WDataOut_1;

// Connect child module input to parent module output 

assign t5_O1_4_WDataIn_1 = Token0_2_WDataOut_1;
endmodule

module DSE_Solution_L2( 
clk,
rst,
DSE_Solution_L2_t5_In0_1,
DSE_Solution_L2_t3_O0_3
); 

input clk;
input rst;
input [31:0] DSE_Solution_L2_t5_In0_1; 
output [31:0] DSE_Solution_L2_t3_O0_3; 
wire [31:0] t5_In0_1_WDataIn_1;
assign t5_In0_1_WDataIn_1 = DSE_Solution_L2_t5_In0_1;
defparam t5_In0_1.DataIn_1_BW = 32;
wire [31:0] t5_In0_1_WDataOut_1;
defparam t5_In0_1.DataOut_1_BW = 32;
HA_INW t5_In0_1 (
	.DataIn_1(t5_In0_1_WDataIn_1) ,
	.DataOut_1(t5_In0_1_WDataOut_1) 
);
wire [31:0] Token0_2_WDataIn_1;
defparam Token0_2.DataIn_1_BW = 32;
wire [31:0] Token0_2_WDataOut_1;
defparam Token0_2.DataOut_1_BW = 32;
HA_TW Token0_2 (
	.DataIn_1(Token0_2_WDataIn_1) ,
	.DataOut_1(Token0_2_WDataOut_1) 
);
wire [31:0] t3_O0_3_WDataIn_1;
defparam t3_O0_3.DataIn_1_BW = 32;
wire [31:0] t3_O0_3_WDataOut_1;
assign DSE_Solution_L2_t3_O0_3 = t3_O0_3_WDataOut_1;
defparam t3_O0_3.DataOut_1_BW = 32;
HA_OW t3_O0_3 (
	.DataIn_1(t3_O0_3_WDataIn_1) ,
	.DataOut_1(t3_O0_3_WDataOut_1) 
);

// Connect child module input to parent module output 

assign Token0_2_WDataIn_1 = t5_In0_1_WDataOut_1;

// Connect child module input to parent module output 

assign t3_O0_3_WDataIn_1 = Token0_2_WDataOut_1;
endmodule

module DSE_Solution_L3( 
clk,
rst,
DSE_Solution_L3_t5_In0_1,
DSE_Solution_L3_t5_O0_3
); 

input clk;
input rst;
input [31:0] DSE_Solution_L3_t5_In0_1; 
output [31:0] DSE_Solution_L3_t5_O0_3; 
wire [31:0] t5_In0_1_WDataIn_1;
assign t5_In0_1_WDataIn_1 = DSE_Solution_L3_t5_In0_1;
defparam t5_In0_1.DataIn_1_BW = 32;
wire [31:0] t5_In0_1_WDataOut_1;
defparam t5_In0_1.DataOut_1_BW = 32;
HA_INW t5_In0_1 (
	.DataIn_1(t5_In0_1_WDataIn_1) ,
	.DataOut_1(t5_In0_1_WDataOut_1) 
);
wire [31:0] Token0_2_WDataIn_1;
defparam Token0_2.DataIn_1_BW = 32;
wire [31:0] Token0_2_WDataOut_1;
defparam Token0_2.DataOut_1_BW = 32;
HA_TW Token0_2 (
	.DataIn_1(Token0_2_WDataIn_1) ,
	.DataOut_1(Token0_2_WDataOut_1) 
);
wire [31:0] t5_O0_3_WDataIn_1;
defparam t5_O0_3.DataIn_1_BW = 32;
wire [31:0] t5_O0_3_WDataOut_1;
assign DSE_Solution_L3_t5_O0_3 = t5_O0_3_WDataOut_1;
defparam t5_O0_3.DataOut_1_BW = 32;
HA_OW t5_O0_3 (
	.DataIn_1(t5_O0_3_WDataIn_1) ,
	.DataOut_1(t5_O0_3_WDataOut_1) 
);

// Connect child module input to parent module output 

assign Token0_2_WDataIn_1 = t5_In0_1_WDataOut_1;

// Connect child module input to parent module output 

assign t5_O0_3_WDataIn_1 = Token0_2_WDataOut_1;
endmodule

module DSE_Solution_L4( 
clk,
rst,
DSE_Solution_L4_t5_In0_1,
DSE_Solution_L4_t5_O0_3
); 

input clk;
input rst;
input [31:0] DSE_Solution_L4_t5_In0_1; 
output [31:0] DSE_Solution_L4_t5_O0_3; 
wire [31:0] t5_In0_1_WDataIn_1;
assign t5_In0_1_WDataIn_1 = DSE_Solution_L4_t5_In0_1;
defparam t5_In0_1.DataIn_1_BW = 32;
wire [31:0] t5_In0_1_WDataOut_1;
defparam t5_In0_1.DataOut_1_BW = 32;
HA_INW t5_In0_1 (
	.DataIn_1(t5_In0_1_WDataIn_1) ,
	.DataOut_1(t5_In0_1_WDataOut_1) 
);
wire [31:0] Token0_2_WDataIn_1;
defparam Token0_2.DataIn_1_BW = 32;
wire [31:0] Token0_2_WDataOut_1;
defparam Token0_2.DataOut_1_BW = 32;
HA_TW Token0_2 (
	.DataIn_1(Token0_2_WDataIn_1) ,
	.DataOut_1(Token0_2_WDataOut_1) 
);
wire [31:0] t5_O0_3_WDataIn_1;
defparam t5_O0_3.DataIn_1_BW = 32;
wire [31:0] t5_O0_3_WDataOut_1;
assign DSE_Solution_L4_t5_O0_3 = t5_O0_3_WDataOut_1;
defparam t5_O0_3.DataOut_1_BW = 32;
HA_OW t5_O0_3 (
	.DataIn_1(t5_O0_3_WDataIn_1) ,
	.DataOut_1(t5_O0_3_WDataOut_1) 
);

// Connect child module input to parent module output 

assign Token0_2_WDataIn_1 = t5_In0_1_WDataOut_1;

// Connect child module input to parent module output 

assign t5_O0_3_WDataIn_1 = Token0_2_WDataOut_1;
endmodule

module DSE_Solution_L5( 
clk,
rst,
DSE_Solution_L5_t5_In0_1,
DSE_Solution_L5_t5_O0_3
); 

input clk;
input rst;
input [31:0] DSE_Solution_L5_t5_In0_1; 
output [31:0] DSE_Solution_L5_t5_O0_3; 
wire [31:0] t5_In0_1_WDataIn_1;
assign t5_In0_1_WDataIn_1 = DSE_Solution_L5_t5_In0_1;
defparam t5_In0_1.DataIn_1_BW = 32;
wire [31:0] t5_In0_1_WDataOut_1;
defparam t5_In0_1.DataOut_1_BW = 32;
HA_INW t5_In0_1 (
	.DataIn_1(t5_In0_1_WDataIn_1) ,
	.DataOut_1(t5_In0_1_WDataOut_1) 
);
wire [31:0] Token0_2_WDataIn_1;
defparam Token0_2.DataIn_1_BW = 32;
wire [31:0] Token0_2_WDataOut_1;
defparam Token0_2.DataOut_1_BW = 32;
HA_TW Token0_2 (
	.DataIn_1(Token0_2_WDataIn_1) ,
	.DataOut_1(Token0_2_WDataOut_1) 
);
wire [31:0] t5_O0_3_WDataIn_1;
defparam t5_O0_3.DataIn_1_BW = 32;
wire [31:0] t5_O0_3_WDataOut_1;
assign DSE_Solution_L5_t5_O0_3 = t5_O0_3_WDataOut_1;
defparam t5_O0_3.DataOut_1_BW = 32;
HA_OW t5_O0_3 (
	.DataIn_1(t5_O0_3_WDataIn_1) ,
	.DataOut_1(t5_O0_3_WDataOut_1) 
);

// Connect child module input to parent module output 

assign Token0_2_WDataIn_1 = t5_In0_1_WDataOut_1;

// Connect child module input to parent module output 

assign t5_O0_3_WDataIn_1 = Token0_2_WDataOut_1;
endmodule

